VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1426.380 2924.800 1427.580 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3486.100 2.400 3487.300 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3224.980 2.400 3226.180 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2964.540 2.400 2965.740 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1692.260 2924.800 1693.460 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2703.420 2.400 2704.620 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2442.980 2.400 2444.180 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2182.540 2.400 2183.740 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1921.420 2.400 1922.620 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1660.980 2.400 1662.180 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1399.860 2.400 1401.060 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1139.420 2.400 1140.620 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 878.980 2.400 880.180 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 617.860 2.400 619.060 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1958.140 2924.800 1959.340 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2223.340 2924.800 2224.540 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2489.220 2924.800 2490.420 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2755.100 2924.800 2756.300 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3020.300 2924.800 3021.500 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3286.180 2924.800 3287.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 32.380 2924.800 33.580 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2289.980 2924.800 2291.180 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2555.860 2924.800 2557.060 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2821.060 2924.800 2822.260 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3086.940 2924.800 3088.140 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3352.820 2924.800 3354.020 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 230.940 2924.800 232.140 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3420.820 2.400 3422.020 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3159.700 2.400 3160.900 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2899.260 2.400 2900.460 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2638.820 2.400 2640.020 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2377.700 2.400 2378.900 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2117.260 2.400 2118.460 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 430.180 2924.800 431.380 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1856.140 2.400 1857.340 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1595.700 2.400 1596.900 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1335.260 2.400 1336.460 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1074.140 2.400 1075.340 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 813.700 2.400 814.900 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 552.580 2.400 553.780 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 357.420 2.400 358.620 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 161.580 2.400 162.780 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 629.420 2924.800 630.620 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 828.660 2924.800 829.860 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1027.900 2924.800 1029.100 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1227.140 2924.800 1228.340 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1493.020 2924.800 1494.220 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1758.900 2924.800 1760.100 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2024.100 2924.800 2025.300 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 164.980 2924.800 166.180 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2422.580 2924.800 2423.780 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2688.460 2924.800 2689.660 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2954.340 2924.800 2955.540 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3219.540 2924.800 3220.740 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3485.420 2924.800 3486.620 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 364.220 2924.800 365.420 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3290.260 2.400 3291.460 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3029.820 2.400 3031.020 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2768.700 2.400 2769.900 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2508.260 2.400 2509.460 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2247.140 2.400 2248.340 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1986.700 2.400 1987.900 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 563.460 2924.800 564.660 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1726.260 2.400 1727.460 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1465.140 2.400 1466.340 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1204.700 2.400 1205.900 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 943.580 2.400 944.780 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 683.140 2.400 684.340 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 422.700 2.400 423.900 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 226.860 2.400 228.060 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 31.700 2.400 32.900 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 762.700 2924.800 763.900 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 961.940 2924.800 963.140 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1161.180 2924.800 1162.380 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1360.420 2924.800 1361.620 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1625.620 2924.800 1626.820 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1891.500 2924.800 1892.700 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2157.380 2924.800 2158.580 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 98.340 2924.800 99.540 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2356.620 2924.800 2357.820 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2621.820 2924.800 2623.020 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2887.700 2924.800 2888.900 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3153.580 2924.800 3154.780 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3418.780 2924.800 3419.980 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 297.580 2924.800 298.780 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3355.540 2.400 3356.740 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3095.100 2.400 3096.300 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2833.980 2.400 2835.180 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2573.540 2.400 2574.740 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2312.420 2.400 2313.620 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2051.980 2.400 2053.180 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 496.820 2924.800 498.020 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1791.540 2.400 1792.740 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1530.420 2.400 1531.620 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1269.980 2.400 1271.180 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1008.860 2.400 1010.060 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 748.420 2.400 749.620 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 487.300 2.400 488.500 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 292.140 2.400 293.340 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 96.300 2.400 97.500 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 696.060 2924.800 697.260 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 895.300 2924.800 896.500 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1094.540 2924.800 1095.740 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1293.780 2924.800 1294.980 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1559.660 2924.800 1560.860 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1824.860 2924.800 1826.060 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2090.740 2924.800 2091.940 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.230 -4.800 629.790 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2402.530 -4.800 2403.090 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2420.010 -4.800 2420.570 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2437.950 -4.800 2438.510 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2455.430 -4.800 2455.990 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.370 -4.800 2473.930 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2490.850 -4.800 2491.410 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2508.790 -4.800 2509.350 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2526.730 -4.800 2527.290 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2544.210 -4.800 2544.770 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2562.150 -4.800 2562.710 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.330 -4.800 806.890 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2579.630 -4.800 2580.190 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2597.570 -4.800 2598.130 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2615.050 -4.800 2615.610 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2632.990 -4.800 2633.550 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2650.470 -4.800 2651.030 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2668.410 -4.800 2668.970 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2685.890 -4.800 2686.450 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2703.830 -4.800 2704.390 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2721.770 -4.800 2722.330 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2739.250 -4.800 2739.810 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.270 -4.800 824.830 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2757.190 -4.800 2757.750 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2774.670 -4.800 2775.230 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2792.610 -4.800 2793.170 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2810.090 -4.800 2810.650 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2828.030 -4.800 2828.590 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2845.510 -4.800 2846.070 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2863.450 -4.800 2864.010 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2881.390 -4.800 2881.950 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.750 -4.800 842.310 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.690 -4.800 860.250 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.170 -4.800 877.730 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.110 -4.800 895.670 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.530 -4.800 931.090 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.470 -4.800 949.030 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.710 -4.800 647.270 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.370 -4.800 1001.930 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.790 -4.800 1037.350 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.730 -4.800 1055.290 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.210 -4.800 1072.770 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.150 -4.800 1090.710 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.630 -4.800 1108.190 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.570 -4.800 1126.130 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.510 -4.800 1144.070 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.650 -4.800 665.210 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.990 -4.800 1161.550 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.930 -4.800 1179.490 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.410 -4.800 1196.970 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.350 -4.800 1214.910 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.830 -4.800 1232.390 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.770 -4.800 1250.330 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1267.250 -4.800 1267.810 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.190 -4.800 1285.750 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1303.130 -4.800 1303.690 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.610 -4.800 1321.170 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.130 -4.800 682.690 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.550 -4.800 1339.110 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.030 -4.800 1356.590 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.970 -4.800 1374.530 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.450 -4.800 1392.010 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.390 -4.800 1409.950 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.870 -4.800 1427.430 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.810 -4.800 1445.370 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.750 -4.800 1463.310 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1480.230 -4.800 1480.790 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1498.170 -4.800 1498.730 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.070 -4.800 700.630 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1515.650 -4.800 1516.210 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1533.590 -4.800 1534.150 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1551.070 -4.800 1551.630 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1569.010 -4.800 1569.570 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1586.490 -4.800 1587.050 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1604.430 -4.800 1604.990 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1621.910 -4.800 1622.470 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.850 -4.800 1640.410 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.790 -4.800 1658.350 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.270 -4.800 1675.830 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.550 -4.800 718.110 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.210 -4.800 1693.770 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1710.690 -4.800 1711.250 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.630 -4.800 1729.190 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1746.110 -4.800 1746.670 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.050 -4.800 1764.610 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1781.530 -4.800 1782.090 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1799.470 -4.800 1800.030 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1817.410 -4.800 1817.970 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1834.890 -4.800 1835.450 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1852.830 -4.800 1853.390 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.490 -4.800 736.050 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.310 -4.800 1870.870 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1888.250 -4.800 1888.810 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.670 -4.800 1924.230 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1976.570 -4.800 1977.130 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.510 -4.800 1995.070 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2029.930 -4.800 2030.490 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.970 -4.800 753.530 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2047.870 -4.800 2048.430 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2065.350 -4.800 2065.910 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2083.290 -4.800 2083.850 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2100.770 -4.800 2101.330 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2118.710 -4.800 2119.270 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2136.190 -4.800 2136.750 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2154.130 -4.800 2154.690 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2172.070 -4.800 2172.630 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2189.550 -4.800 2190.110 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2207.490 -4.800 2208.050 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.910 -4.800 771.470 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2224.970 -4.800 2225.530 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2242.910 -4.800 2243.470 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2260.390 -4.800 2260.950 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2278.330 -4.800 2278.890 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2295.810 -4.800 2296.370 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2313.750 -4.800 2314.310 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2331.230 -4.800 2331.790 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2349.170 -4.800 2349.730 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2367.110 -4.800 2367.670 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2384.590 -4.800 2385.150 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.850 -4.800 789.410 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.750 -4.800 635.310 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2408.510 -4.800 2409.070 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2425.990 -4.800 2426.550 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2443.930 -4.800 2444.490 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2461.410 -4.800 2461.970 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2479.350 -4.800 2479.910 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2496.830 -4.800 2497.390 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2514.770 -4.800 2515.330 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2532.250 -4.800 2532.810 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2550.190 -4.800 2550.750 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2567.670 -4.800 2568.230 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.310 -4.800 812.870 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2585.610 -4.800 2586.170 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2603.550 -4.800 2604.110 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2621.030 -4.800 2621.590 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2638.970 -4.800 2639.530 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2656.450 -4.800 2657.010 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2674.390 -4.800 2674.950 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2691.870 -4.800 2692.430 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2709.810 -4.800 2710.370 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2727.290 -4.800 2727.850 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2745.230 -4.800 2745.790 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.250 -4.800 830.810 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2763.170 -4.800 2763.730 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2780.650 -4.800 2781.210 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.590 -4.800 2799.150 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2816.070 -4.800 2816.630 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2834.010 -4.800 2834.570 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2851.490 -4.800 2852.050 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2869.430 -4.800 2869.990 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.730 -4.800 848.290 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.670 -4.800 866.230 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.150 -4.800 883.710 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.090 -4.800 901.650 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.510 -4.800 937.070 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.690 -4.800 653.250 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.410 -4.800 989.970 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.770 -4.800 1043.330 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.710 -4.800 1061.270 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.190 -4.800 1078.750 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.130 -4.800 1096.690 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.610 -4.800 1114.170 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.550 -4.800 1132.110 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.030 -4.800 1149.590 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.630 -4.800 671.190 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.970 -4.800 1167.530 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.910 -4.800 1185.470 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.390 -4.800 1202.950 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.330 -4.800 1220.890 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.810 -4.800 1238.370 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.750 -4.800 1256.310 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.230 -4.800 1273.790 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.170 -4.800 1291.730 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1308.650 -4.800 1309.210 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.590 -4.800 1327.150 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.110 -4.800 688.670 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.070 -4.800 1344.630 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.010 -4.800 1362.570 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.950 -4.800 1380.510 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.430 -4.800 1397.990 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.370 -4.800 1415.930 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.850 -4.800 1433.410 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1450.790 -4.800 1451.350 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.270 -4.800 1468.830 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1486.210 -4.800 1486.770 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.690 -4.800 1504.250 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.050 -4.800 706.610 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.630 -4.800 1522.190 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.570 -4.800 1540.130 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.050 -4.800 1557.610 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.990 -4.800 1575.550 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1592.470 -4.800 1593.030 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.410 -4.800 1610.970 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.890 -4.800 1628.450 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.830 -4.800 1646.390 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1663.310 -4.800 1663.870 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1681.250 -4.800 1681.810 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.530 -4.800 724.090 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1699.190 -4.800 1699.750 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.670 -4.800 1717.230 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1734.610 -4.800 1735.170 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1752.090 -4.800 1752.650 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.030 -4.800 1770.590 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.510 -4.800 1788.070 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1805.450 -4.800 1806.010 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.930 -4.800 1823.490 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1840.870 -4.800 1841.430 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1858.350 -4.800 1858.910 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.470 -4.800 742.030 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1876.290 -4.800 1876.850 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1894.230 -4.800 1894.790 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1929.650 -4.800 1930.210 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1982.550 -4.800 1983.110 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2000.490 -4.800 2001.050 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2017.970 -4.800 2018.530 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2035.910 -4.800 2036.470 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.950 -4.800 759.510 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2053.850 -4.800 2054.410 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2071.330 -4.800 2071.890 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.270 -4.800 2089.830 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2106.750 -4.800 2107.310 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2124.690 -4.800 2125.250 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2142.170 -4.800 2142.730 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2160.110 -4.800 2160.670 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2177.590 -4.800 2178.150 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2195.530 -4.800 2196.090 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2213.010 -4.800 2213.570 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.890 -4.800 777.450 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.950 -4.800 2231.510 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2248.890 -4.800 2249.450 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2266.370 -4.800 2266.930 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2284.310 -4.800 2284.870 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2301.790 -4.800 2302.350 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2319.730 -4.800 2320.290 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2337.210 -4.800 2337.770 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2355.150 -4.800 2355.710 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2372.630 -4.800 2373.190 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2390.570 -4.800 2391.130 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.370 -4.800 794.930 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.730 -4.800 641.290 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2414.030 -4.800 2414.590 2.400 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2431.970 -4.800 2432.530 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2449.450 -4.800 2450.010 2.400 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2467.390 -4.800 2467.950 2.400 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2485.330 -4.800 2485.890 2.400 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2502.810 -4.800 2503.370 2.400 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2520.750 -4.800 2521.310 2.400 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2538.230 -4.800 2538.790 2.400 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2556.170 -4.800 2556.730 2.400 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2573.650 -4.800 2574.210 2.400 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.290 -4.800 818.850 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2591.590 -4.800 2592.150 2.400 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2609.070 -4.800 2609.630 2.400 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2627.010 -4.800 2627.570 2.400 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2644.950 -4.800 2645.510 2.400 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2662.430 -4.800 2662.990 2.400 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2680.370 -4.800 2680.930 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2697.850 -4.800 2698.410 2.400 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2715.790 -4.800 2716.350 2.400 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2733.270 -4.800 2733.830 2.400 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2751.210 -4.800 2751.770 2.400 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.770 -4.800 836.330 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2768.690 -4.800 2769.250 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2786.630 -4.800 2787.190 2.400 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2804.110 -4.800 2804.670 2.400 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2822.050 -4.800 2822.610 2.400 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2839.990 -4.800 2840.550 2.400 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2857.470 -4.800 2858.030 2.400 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2875.410 -4.800 2875.970 2.400 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.710 -4.800 854.270 2.400 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.190 -4.800 871.750 2.400 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.130 -4.800 889.690 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.070 -4.800 907.630 2.400 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.550 -4.800 925.110 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.490 -4.800 943.050 2.400 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.670 -4.800 659.230 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.390 -4.800 995.950 2.400 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.810 -4.800 1031.370 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.750 -4.800 1049.310 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.690 -4.800 1067.250 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.170 -4.800 1084.730 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.110 -4.800 1102.670 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.590 -4.800 1120.150 2.400 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.530 -4.800 1138.090 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.010 -4.800 1155.570 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.150 -4.800 676.710 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.950 -4.800 1173.510 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.430 -4.800 1190.990 2.400 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.370 -4.800 1208.930 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1225.850 -4.800 1226.410 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.790 -4.800 1244.350 2.400 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.730 -4.800 1262.290 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1279.210 -4.800 1279.770 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.150 -4.800 1297.710 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.630 -4.800 1315.190 2.400 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.570 -4.800 1333.130 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.090 -4.800 694.650 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1350.050 -4.800 1350.610 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.990 -4.800 1368.550 2.400 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.470 -4.800 1386.030 2.400 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.410 -4.800 1403.970 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.350 -4.800 1421.910 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.830 -4.800 1439.390 2.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.770 -4.800 1457.330 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.250 -4.800 1474.810 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.190 -4.800 1492.750 2.400 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1509.670 -4.800 1510.230 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.030 -4.800 712.590 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1527.610 -4.800 1528.170 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.090 -4.800 1545.650 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1563.030 -4.800 1563.590 2.400 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.970 -4.800 1581.530 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1598.450 -4.800 1599.010 2.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.390 -4.800 1616.950 2.400 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.870 -4.800 1634.430 2.400 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.810 -4.800 1652.370 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1669.290 -4.800 1669.850 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.230 -4.800 1687.790 2.400 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.510 -4.800 730.070 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.710 -4.800 1705.270 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.650 -4.800 1723.210 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1740.130 -4.800 1740.690 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.070 -4.800 1758.630 2.400 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.010 -4.800 1776.570 2.400 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.490 -4.800 1794.050 2.400 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1811.430 -4.800 1811.990 2.400 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.910 -4.800 1829.470 2.400 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1846.850 -4.800 1847.410 2.400 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.330 -4.800 1864.890 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.450 -4.800 748.010 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1882.270 -4.800 1882.830 2.400 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.630 -4.800 1936.190 2.400 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1988.530 -4.800 1989.090 2.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2023.950 -4.800 2024.510 2.400 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.890 -4.800 2042.450 2.400 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.930 -4.800 765.490 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2059.370 -4.800 2059.930 2.400 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2077.310 -4.800 2077.870 2.400 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2094.790 -4.800 2095.350 2.400 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.730 -4.800 2113.290 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.670 -4.800 2131.230 2.400 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2148.150 -4.800 2148.710 2.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2166.090 -4.800 2166.650 2.400 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.570 -4.800 2184.130 2.400 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2201.510 -4.800 2202.070 2.400 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.990 -4.800 2219.550 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.870 -4.800 783.430 2.400 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2236.930 -4.800 2237.490 2.400 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2254.410 -4.800 2254.970 2.400 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2272.350 -4.800 2272.910 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2290.290 -4.800 2290.850 2.400 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2307.770 -4.800 2308.330 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2325.710 -4.800 2326.270 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2343.190 -4.800 2343.750 2.400 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2361.130 -4.800 2361.690 2.400 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2378.610 -4.800 2379.170 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2396.550 -4.800 2397.110 2.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.350 -4.800 800.910 2.400 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -10.030 -4.670 2929.650 -1.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 14.090 2934.450 17.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 194.090 2934.450 197.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 374.090 2934.450 377.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 554.090 2934.450 557.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 734.090 2934.450 737.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 914.090 2934.450 917.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1094.090 2934.450 1097.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1274.090 2934.450 1277.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1454.090 2934.450 1457.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1634.090 2934.450 1637.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1814.090 2934.450 1817.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1994.090 2934.450 1997.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2174.090 2934.450 2177.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2354.090 2934.450 2357.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2534.090 2934.450 2537.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2714.090 2934.450 2717.190 ;
    END
    PORT
      LAYER met5 ;
        RECT 188.970 2808.790 552.070 2811.890 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2894.090 2934.450 2897.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3074.090 2934.450 3077.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3254.090 2934.450 3257.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3434.090 2934.450 3437.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 3521.250 2929.650 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 -9.470 192.070 167.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 -9.470 372.070 167.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 -9.470 552.070 167.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1628.970 -9.470 1632.070 190.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 -9.470 1812.070 190.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 -9.470 1992.070 190.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 -9.470 2352.070 190.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 -9.470 2532.070 190.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 -9.470 2712.070 190.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 410.180 192.070 567.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 410.180 372.070 567.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 410.180 552.070 567.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 -9.470 732.070 567.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 613.380 1812.070 786.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 613.380 1992.070 786.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 -9.470 2172.070 786.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 613.380 2352.070 786.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 1005.760 192.070 1465.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 1005.760 372.070 1465.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 1005.760 552.070 1465.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 1005.760 732.070 1465.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 -9.470 912.070 1465.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 1224.340 1812.070 1494.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 1224.340 1992.070 1494.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 1224.340 2172.070 1494.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 1840.520 1812.070 2050.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 1840.520 1992.070 2050.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 1840.520 2172.070 2050.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 1224.340 2352.070 2050.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 2156.900 192.070 2310.980 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 2156.900 372.070 2310.980 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 2156.900 552.070 2310.980 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 2734.120 192.070 2885.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 2734.120 372.070 2885.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 2734.120 552.070 2885.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 2742.660 1812.070 3019.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 2742.660 1992.070 3019.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 2742.660 2172.070 3019.180 ;
    END
    PORT
      LAYER met4 ;
        RECT -10.030 -4.670 -6.930 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2926.550 -4.670 2929.650 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.970 -9.470 12.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 3352.140 192.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 3352.140 372.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 3352.140 552.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 2156.900 732.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 2156.900 912.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 -9.470 1092.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 -9.470 1272.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1448.970 -9.470 1452.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1628.970 613.380 1632.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 3364.800 1812.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 3364.800 1992.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 3364.800 2172.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 2742.660 2352.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 613.380 2532.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 613.380 2712.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2888.970 -9.470 2892.070 3529.150 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -19.630 -14.270 2939.250 -11.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 32.930 2944.050 36.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 212.930 2944.050 216.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 392.930 2944.050 396.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 207.570 487.630 570.670 490.730 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 572.930 2944.050 576.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 752.930 2944.050 756.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 932.930 2944.050 936.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1112.930 2944.050 1116.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1292.930 2944.050 1296.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1472.930 2944.050 1476.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1652.930 2944.050 1656.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1832.930 2944.050 1836.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2012.930 2944.050 2016.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2192.930 2944.050 2196.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2372.930 2944.050 2376.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2552.930 2944.050 2556.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2732.930 2944.050 2736.030 ;
    END
    PORT
      LAYER met5 ;
        RECT 207.570 2818.230 570.670 2821.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2912.930 2944.050 2916.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3092.930 2944.050 3096.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3272.930 2944.050 3276.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3452.930 2944.050 3456.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -19.630 3530.850 2939.250 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 207.570 -19.070 210.670 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.570 -19.070 390.670 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 567.570 -19.070 570.670 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1647.570 -19.070 1650.670 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1827.570 -19.070 1830.670 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2007.570 -19.070 2010.670 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2367.570 -19.070 2370.670 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.570 -19.070 2550.670 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2727.570 -19.070 2730.670 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 207.570 410.420 210.670 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.570 410.420 390.670 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 567.570 410.420 570.670 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 747.570 -19.070 750.670 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1827.570 613.620 1830.670 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2007.570 613.620 2010.670 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2187.570 -19.070 2190.670 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2367.570 613.620 2370.670 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 207.570 1006.000 210.670 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.570 1006.000 390.670 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 567.570 1006.000 570.670 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 747.570 1006.000 750.670 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1827.570 1224.580 1830.670 1494.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 2007.570 1224.580 2010.670 1494.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 2187.570 1224.580 2190.670 1494.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 1827.570 1840.760 1830.670 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2007.570 1840.760 2010.670 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2187.570 1840.760 2190.670 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2367.570 1224.580 2370.670 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 207.570 2157.140 210.670 2310.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.570 2157.140 390.670 2310.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 567.570 2157.140 570.670 2310.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 207.570 2734.360 210.670 2885.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.570 2734.360 390.670 2885.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 567.570 2734.360 570.670 2885.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1827.570 2742.900 1830.670 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2007.570 2742.900 2010.670 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2187.570 2742.900 2190.670 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT -19.630 -14.270 -16.530 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2936.150 -14.270 2939.250 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 27.570 -19.070 30.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 207.570 3352.380 210.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.570 3352.380 390.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 567.570 3352.380 570.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 747.570 2157.140 750.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 927.570 -19.070 930.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1107.570 -19.070 1110.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1287.570 -19.070 1290.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1467.570 -19.070 1470.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1647.570 613.620 1650.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1827.570 3365.040 1830.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2007.570 3365.040 2010.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2187.570 3365.040 2190.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2367.570 2742.900 2370.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2547.570 613.620 2550.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2727.570 613.620 2730.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2907.570 -19.070 2910.670 3538.750 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -29.230 -23.870 2948.850 -20.770 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 51.530 2953.650 54.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 231.530 2953.650 234.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 411.530 2953.650 414.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 591.530 2953.650 594.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 771.530 2953.650 774.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 951.530 2953.650 954.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1131.530 2953.650 1134.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1311.530 2953.650 1314.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1491.530 2953.650 1494.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1671.530 2953.650 1674.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1851.530 2953.650 1854.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2031.530 2953.650 2034.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2211.530 2953.650 2214.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2391.530 2953.650 2394.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2571.530 2953.650 2574.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2751.530 2953.650 2754.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2931.530 2953.650 2934.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3111.530 2953.650 3114.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3291.530 2953.650 3294.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3471.530 2953.650 3474.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -29.230 3540.450 2948.850 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 226.170 -28.670 229.270 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 406.170 -28.670 409.270 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 586.170 -28.670 589.270 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1666.170 -28.670 1669.270 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1846.170 -28.670 1849.270 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2026.170 -28.670 2029.270 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2386.170 -28.670 2389.270 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2566.170 -28.670 2569.270 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2746.170 -28.670 2749.270 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 226.170 410.420 229.270 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 406.170 410.420 409.270 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 586.170 410.420 589.270 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 766.170 -28.670 769.270 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1846.170 613.620 1849.270 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2026.170 613.620 2029.270 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2206.170 -28.670 2209.270 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2386.170 613.620 2389.270 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 226.170 1006.000 229.270 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 406.170 1006.000 409.270 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 586.170 1006.000 589.270 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 766.170 1006.000 769.270 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1846.170 1224.580 1849.270 1494.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 2026.170 1224.580 2029.270 1494.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 1846.170 1840.760 1849.270 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2026.170 1840.760 2029.270 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2206.170 1224.580 2209.270 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2386.170 1224.580 2389.270 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 226.170 2157.140 229.270 2310.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 406.170 2157.140 409.270 2310.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 586.170 2157.140 589.270 2310.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 226.170 2734.360 229.270 2885.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 406.170 2734.360 409.270 2885.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 586.170 2734.360 589.270 2885.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1846.170 2742.900 1849.270 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2026.170 2742.900 2029.270 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT -29.230 -23.870 -26.130 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 2945.750 -23.870 2948.850 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 46.170 -28.670 49.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 226.170 3352.380 229.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 406.170 3352.380 409.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 586.170 3352.380 589.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 766.170 2157.140 769.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 946.170 -28.670 949.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1126.170 -28.670 1129.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1306.170 -28.670 1309.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1486.170 -28.670 1489.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1666.170 613.620 1669.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1846.170 3365.040 1849.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2026.170 3365.040 2029.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2206.170 2742.900 2209.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2386.170 2742.900 2389.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2566.170 613.620 2569.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2746.170 613.620 2749.270 3548.350 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -38.830 -33.470 2958.450 -30.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 70.130 2963.250 73.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 250.130 2963.250 253.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 430.130 2963.250 433.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 610.130 2963.250 613.230 ;
    END
    PORT
      LAYER met5 ;
        RECT 1864.770 695.430 2407.870 698.530 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 790.130 2963.250 793.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 970.130 2963.250 973.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1150.130 2963.250 1153.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1330.130 2963.250 1333.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1510.130 2963.250 1513.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1690.130 2963.250 1693.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1870.130 2963.250 1873.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2050.130 2963.250 2053.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2230.130 2963.250 2233.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2410.130 2963.250 2413.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2590.130 2963.250 2593.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2770.130 2963.250 2773.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2950.130 2963.250 2953.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3130.130 2963.250 3133.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3310.130 2963.250 3313.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3490.130 2963.250 3493.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -38.830 3550.050 2958.450 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 244.770 -38.270 247.870 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.770 -38.270 427.870 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.770 -38.270 607.870 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1684.770 -38.270 1687.870 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.770 -38.270 1867.870 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2044.770 -38.270 2047.870 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2404.770 -38.270 2407.870 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2584.770 -38.270 2587.870 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2764.770 -38.270 2767.870 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 244.770 410.420 247.870 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.770 410.420 427.870 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.770 410.420 607.870 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 784.770 -38.270 787.870 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.770 613.620 1867.870 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2044.770 613.620 2047.870 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2224.770 -38.270 2227.870 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2404.770 613.620 2407.870 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 244.770 1006.000 247.870 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.770 1006.000 427.870 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.770 1006.000 607.870 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 784.770 1006.000 787.870 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.770 1224.580 1867.870 1494.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 2044.770 1224.580 2047.870 1494.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.770 1840.760 1867.870 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2044.770 1840.760 2047.870 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2224.770 1224.580 2227.870 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2404.770 1224.580 2407.870 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 244.770 2157.140 247.870 2310.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.770 2157.140 427.870 2310.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.770 2157.140 607.870 2310.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 244.770 2734.360 247.870 2885.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.770 2734.360 427.870 2885.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.770 2734.360 607.870 2885.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.770 2742.900 1867.870 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2044.770 2742.900 2047.870 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT -38.830 -33.470 -35.730 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2955.350 -33.470 2958.450 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.770 -38.270 67.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 244.770 3352.380 247.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.770 3352.380 427.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.770 3352.380 607.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 784.770 2157.140 787.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 964.770 -38.270 967.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1144.770 -38.270 1147.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1324.770 -38.270 1327.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1504.770 -38.270 1507.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1684.770 613.620 1687.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.770 3365.040 1867.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2044.770 3365.040 2047.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2224.770 2742.900 2227.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2404.770 2742.900 2407.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2584.770 613.620 2587.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2764.770 613.620 2767.870 3557.950 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -34.030 -28.670 2953.650 -25.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 141.530 2953.650 144.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 321.530 2953.650 324.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 501.530 2953.650 504.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 681.530 2953.650 684.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 861.530 2953.650 864.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1041.530 2953.650 1044.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1221.530 2953.650 1224.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1401.530 2953.650 1404.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1581.530 2953.650 1584.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1761.530 2953.650 1764.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 1941.530 2953.650 1944.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2121.530 2953.650 2124.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2301.530 2953.650 2304.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2481.530 2953.650 2484.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2661.530 2953.650 2664.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 2841.530 2953.650 2844.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3021.530 2953.650 3024.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3201.530 2953.650 3204.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3381.530 2953.650 3384.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3545.250 2953.650 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 316.170 -28.670 319.270 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.170 -28.670 499.270 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 676.170 -28.670 679.270 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1756.170 -28.670 1759.270 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.170 -28.670 1939.270 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2296.170 -28.670 2299.270 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2476.170 -28.670 2479.270 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2656.170 -28.670 2659.270 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 316.170 410.420 319.270 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.170 410.420 499.270 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 676.170 410.420 679.270 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 856.170 -28.670 859.270 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1756.170 613.620 1759.270 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.170 613.620 1939.270 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2116.170 -28.670 2119.270 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2296.170 613.620 2299.270 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 316.170 1006.000 319.270 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.170 1006.000 499.270 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 676.170 1006.000 679.270 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 856.170 1006.000 859.270 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1756.170 1224.580 1759.270 1494.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.170 1224.580 1939.270 1494.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 2116.170 1224.580 2119.270 1494.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 1756.170 1840.760 1759.270 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.170 1840.760 1939.270 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2116.170 1840.760 2119.270 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2296.170 1224.580 2299.270 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 316.170 2157.140 319.270 2310.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.170 2157.140 499.270 2310.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 676.170 2157.140 679.270 2310.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 316.170 2734.360 319.270 2885.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.170 2734.360 499.270 2885.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1756.170 2742.900 1759.270 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.170 2742.900 1939.270 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2116.170 2742.900 2119.270 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT -34.030 -28.670 -30.930 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 136.170 -28.670 139.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 316.170 3352.380 319.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 496.170 3352.380 499.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 676.170 2734.360 679.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 856.170 2157.140 859.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1036.170 -28.670 1039.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1216.170 -28.670 1219.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1396.170 -28.670 1399.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1576.170 -28.670 1579.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1756.170 3365.040 1759.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.170 3365.040 1939.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2116.170 3365.040 2119.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2296.170 2742.900 2299.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2476.170 613.620 2479.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2656.170 613.620 2659.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2836.170 -28.670 2839.270 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2950.550 -28.670 2953.650 3548.350 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -43.630 -38.270 2963.250 -35.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 160.130 2963.250 163.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 340.130 2963.250 343.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 520.130 2963.250 523.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 700.130 2963.250 703.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 880.130 2963.250 883.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1060.130 2963.250 1063.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1240.130 2963.250 1243.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1420.130 2963.250 1423.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1600.130 2963.250 1603.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1780.130 2963.250 1783.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1960.130 2963.250 1963.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2140.130 2963.250 2143.230 ;
    END
    PORT
      LAYER met5 ;
        RECT 334.770 2234.830 697.870 2237.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2320.130 2963.250 2323.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2500.130 2963.250 2503.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2680.130 2963.250 2683.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2860.130 2963.250 2863.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3040.130 2963.250 3043.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3220.130 2963.250 3223.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3400.130 2963.250 3403.230 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3554.850 2963.250 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.770 -38.270 337.870 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 514.770 -38.270 517.870 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1594.770 -38.270 1597.870 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1774.770 -38.270 1777.870 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.770 -38.270 1957.870 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2314.770 -38.270 2317.870 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2494.770 -38.270 2497.870 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2674.770 -38.270 2677.870 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.770 410.420 337.870 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 514.770 410.420 517.870 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 694.770 -38.270 697.870 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 874.770 -38.270 877.870 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1774.770 613.620 1777.870 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.770 613.620 1957.870 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2134.770 -38.270 2137.870 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2314.770 613.620 2317.870 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.770 1006.000 337.870 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 514.770 1006.000 517.870 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 694.770 1006.000 697.870 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 874.770 1006.000 877.870 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1774.770 1224.580 1777.870 1494.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.770 1224.580 1957.870 1494.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 2134.770 1224.580 2137.870 1494.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 1774.770 1840.760 1777.870 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.770 1840.760 1957.870 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2134.770 1840.760 2137.870 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2314.770 1224.580 2317.870 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.770 2157.140 337.870 2310.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 514.770 2157.140 517.870 2310.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 694.770 2157.140 697.870 2310.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.770 2734.360 337.870 2885.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 514.770 2734.360 517.870 2885.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1774.770 2742.900 1777.870 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.770 2742.900 1957.870 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2134.770 2742.900 2137.870 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT -43.630 -38.270 -40.530 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 154.770 -38.270 157.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.770 3352.380 337.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 514.770 3352.380 517.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 694.770 2734.360 697.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 874.770 2157.140 877.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1054.770 -38.270 1057.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1234.770 -38.270 1237.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1414.770 -38.270 1417.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1594.770 613.620 1597.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1774.770 3365.040 1777.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.770 3365.040 1957.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2134.770 3365.040 2137.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2314.770 2742.900 2317.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2494.770 613.620 2497.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2674.770 613.620 2677.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2854.770 -38.270 2857.870 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2960.150 -38.270 2963.250 3557.950 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.830 -9.470 2934.450 -6.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 104.090 2934.450 107.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 284.090 2934.450 287.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 464.090 2934.450 467.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 644.090 2934.450 647.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 824.090 2934.450 827.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1004.090 2934.450 1007.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1184.090 2934.450 1187.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1364.090 2934.450 1367.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1544.090 2934.450 1547.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1724.090 2934.450 1727.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 1904.090 2934.450 1907.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2084.090 2934.450 2087.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2264.090 2934.450 2267.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2444.090 2934.450 2447.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2624.090 2934.450 2627.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2804.090 2934.450 2807.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 2984.090 2934.450 2987.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3164.090 2934.450 3167.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3344.090 2934.450 3347.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3526.050 2934.450 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 -9.470 282.070 167.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 -9.470 462.070 167.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 -9.470 642.070 167.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 -9.470 1722.070 190.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 -9.470 1902.070 190.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.970 -9.470 2082.070 190.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 -9.470 2442.070 190.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 -9.470 2622.070 190.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 410.180 282.070 567.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 410.180 462.070 567.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 410.180 642.070 567.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 818.970 -9.470 822.070 567.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 613.380 1722.070 786.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 613.380 1902.070 786.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.970 613.380 2082.070 786.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 -9.470 2262.070 786.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 1005.760 282.070 1465.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 1005.760 462.070 1465.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 1005.760 642.070 1465.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 818.970 1005.760 822.070 1465.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 1224.340 1722.070 1494.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 1224.340 1902.070 1494.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.970 1224.340 2082.070 1494.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 1840.520 1722.070 2050.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 1840.520 1902.070 2050.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.970 1840.520 2082.070 2050.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 1224.340 2262.070 2050.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 2156.900 282.070 2310.980 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 2156.900 462.070 2310.980 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 2156.900 642.070 2310.980 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 2734.120 282.070 2885.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 2734.120 462.070 2885.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 2734.120 642.070 2885.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 2742.660 1722.070 3019.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 2742.660 1902.070 3019.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.970 2742.660 2082.070 3019.180 ;
    END
    PORT
      LAYER met4 ;
        RECT -14.830 -9.470 -11.730 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.970 -9.470 102.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 3352.140 282.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 3352.140 462.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 3352.140 642.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 818.970 2156.900 822.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 998.970 -9.470 1002.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1178.970 -9.470 1182.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.970 -9.470 1362.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1538.970 -9.470 1542.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 3364.800 1722.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 3364.800 1902.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.970 3364.800 2082.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 2742.660 2262.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 613.380 2442.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 613.380 2622.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2798.970 -9.470 2802.070 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2931.350 -9.470 2934.450 3529.150 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.430 -19.070 2944.050 -15.970 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 122.930 2944.050 126.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 302.930 2944.050 306.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 482.930 2944.050 486.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 662.930 2944.050 666.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 842.930 2944.050 846.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1022.930 2944.050 1026.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1202.930 2944.050 1206.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1382.930 2944.050 1386.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1562.930 2944.050 1566.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1742.930 2944.050 1746.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 1922.930 2944.050 1926.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2102.930 2944.050 2106.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2282.930 2944.050 2286.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2462.930 2944.050 2466.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2642.930 2944.050 2646.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 2822.930 2944.050 2826.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3002.930 2944.050 3006.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3182.930 2944.050 3186.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3362.930 2944.050 3366.030 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3535.650 2944.050 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 297.570 -19.070 300.670 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.570 -19.070 480.670 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 657.570 -19.070 660.670 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1737.570 -19.070 1740.670 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.570 -19.070 1920.670 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2097.570 -19.070 2100.670 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2277.570 -19.070 2280.670 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2457.570 -19.070 2460.670 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2637.570 -19.070 2640.670 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 297.570 410.420 300.670 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.570 410.420 480.670 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 657.570 410.420 660.670 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 837.570 -19.070 840.670 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 1737.570 613.620 1740.670 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.570 613.620 1920.670 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2097.570 613.620 2100.670 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2277.570 613.620 2280.670 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 297.570 1006.000 300.670 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.570 1006.000 480.670 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 657.570 1006.000 660.670 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 837.570 1006.000 840.670 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 1737.570 1224.580 1740.670 1494.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.570 1224.580 1920.670 1494.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 2097.570 1224.580 2100.670 1494.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 1737.570 1840.760 1740.670 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.570 1840.760 1920.670 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2097.570 1840.760 2100.670 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2277.570 1224.580 2280.670 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 297.570 2157.140 300.670 2310.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.570 2157.140 480.670 2310.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 657.570 2157.140 660.670 2310.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 297.570 2734.360 300.670 2885.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.570 2734.360 480.670 2885.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 657.570 2734.360 660.670 2885.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1737.570 2742.900 1740.670 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.570 2742.900 1920.670 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2097.570 2742.900 2100.670 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT -24.430 -19.070 -21.330 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 117.570 -19.070 120.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 297.570 3352.380 300.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.570 3352.380 480.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 657.570 3352.380 660.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 837.570 2157.140 840.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1017.570 -19.070 1020.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1197.570 -19.070 1200.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.570 -19.070 1380.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.570 -19.070 1560.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1737.570 3365.040 1740.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 1917.570 3365.040 1920.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2097.570 3365.040 2100.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2277.570 2742.900 2280.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2457.570 613.620 2460.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2637.570 613.620 2640.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2817.570 -19.070 2820.670 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2940.950 -19.070 2944.050 3538.750 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.150 -4.800 239.710 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.630 -4.800 257.190 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.570 -4.800 275.130 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.050 -4.800 292.610 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.990 -4.800 310.550 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.470 -4.800 328.030 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.410 -4.800 345.970 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.890 -4.800 363.450 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.830 -4.800 381.390 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.310 -4.800 398.870 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.590 -4.800 62.150 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.250 -4.800 416.810 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.190 -4.800 434.750 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.670 -4.800 452.230 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.610 -4.800 470.170 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.090 -4.800 487.650 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.030 -4.800 505.590 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.510 -4.800 523.070 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.450 -4.800 541.010 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.930 -4.800 558.490 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.870 -4.800 576.430 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.050 -4.800 85.610 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.810 -4.800 594.370 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.290 -4.800 611.850 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.970 -4.800 109.530 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.430 -4.800 132.990 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.370 -4.800 150.930 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.850 -4.800 168.410 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.790 -4.800 186.350 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.270 -4.800 203.830 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.210 -4.800 221.770 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.650 -4.800 44.210 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.670 -4.800 245.230 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.610 -4.800 263.170 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.090 -4.800 280.650 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.030 -4.800 298.590 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.970 -4.800 316.530 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.450 -4.800 334.010 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.390 -4.800 351.950 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.870 -4.800 369.430 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.810 -4.800 387.370 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.290 -4.800 404.850 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.570 -4.800 68.130 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.230 -4.800 422.790 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.710 -4.800 440.270 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.650 -4.800 458.210 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.590 -4.800 476.150 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.070 -4.800 493.630 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.010 -4.800 511.570 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.490 -4.800 529.050 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.430 -4.800 546.990 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.910 -4.800 564.470 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.850 -4.800 582.410 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.030 -4.800 91.590 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.330 -4.800 599.890 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.270 -4.800 617.830 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.950 -4.800 115.510 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.410 -4.800 138.970 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.350 -4.800 156.910 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.830 -4.800 174.390 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.770 -4.800 192.330 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.250 -4.800 209.810 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.190 -4.800 227.750 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.630 -4.800 50.190 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.650 -4.800 251.210 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.590 -4.800 269.150 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.070 -4.800 286.630 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.010 -4.800 304.570 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.490 -4.800 322.050 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.430 -4.800 339.990 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.370 -4.800 357.930 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.850 -4.800 375.410 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.790 -4.800 393.350 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.270 -4.800 410.830 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.550 -4.800 74.110 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.210 -4.800 428.770 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 -4.800 446.250 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.630 -4.800 464.190 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.110 -4.800 481.670 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.050 -4.800 499.610 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.530 -4.800 517.090 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.470 -4.800 535.030 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.410 -4.800 552.970 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.890 -4.800 570.450 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.830 -4.800 588.390 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.010 -4.800 97.570 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.310 -4.800 605.870 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.250 -4.800 623.810 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.930 -4.800 121.490 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.390 -4.800 144.950 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.870 -4.800 162.430 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.810 -4.800 180.370 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.750 -4.800 198.310 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.230 -4.800 215.790 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.170 -4.800 233.730 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.610 -4.800 56.170 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.530 -4.800 80.090 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.990 -4.800 103.550 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.450 -4.800 127.010 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2914.100 3508.885 ;
      LAYER met1 ;
        RECT 2.830 1.400 2917.250 3509.040 ;
      LAYER met2 ;
        RECT 2.860 3517.320 40.150 3518.050 ;
        RECT 41.270 3517.320 121.110 3518.050 ;
        RECT 122.230 3517.320 202.070 3518.050 ;
        RECT 203.190 3517.320 283.490 3518.050 ;
        RECT 284.610 3517.320 364.450 3518.050 ;
        RECT 365.570 3517.320 445.410 3518.050 ;
        RECT 446.530 3517.320 526.830 3518.050 ;
        RECT 527.950 3517.320 607.790 3518.050 ;
        RECT 608.910 3517.320 688.750 3518.050 ;
        RECT 689.870 3517.320 770.170 3518.050 ;
        RECT 771.290 3517.320 851.130 3518.050 ;
        RECT 852.250 3517.320 932.090 3518.050 ;
        RECT 933.210 3517.320 1013.510 3518.050 ;
        RECT 1014.630 3517.320 1094.470 3518.050 ;
        RECT 1095.590 3517.320 1175.430 3518.050 ;
        RECT 1176.550 3517.320 1256.850 3518.050 ;
        RECT 1257.970 3517.320 1337.810 3518.050 ;
        RECT 1338.930 3517.320 1418.770 3518.050 ;
        RECT 1419.890 3517.320 1500.190 3518.050 ;
        RECT 1501.310 3517.320 1581.150 3518.050 ;
        RECT 1582.270 3517.320 1662.110 3518.050 ;
        RECT 1663.230 3517.320 1743.530 3518.050 ;
        RECT 1744.650 3517.320 1824.490 3518.050 ;
        RECT 1825.610 3517.320 1905.450 3518.050 ;
        RECT 1906.570 3517.320 1986.870 3518.050 ;
        RECT 1987.990 3517.320 2067.830 3518.050 ;
        RECT 2068.950 3517.320 2148.790 3518.050 ;
        RECT 2149.910 3517.320 2230.210 3518.050 ;
        RECT 2231.330 3517.320 2311.170 3518.050 ;
        RECT 2312.290 3517.320 2392.130 3518.050 ;
        RECT 2393.250 3517.320 2473.550 3518.050 ;
        RECT 2474.670 3517.320 2554.510 3518.050 ;
        RECT 2555.630 3517.320 2635.470 3518.050 ;
        RECT 2636.590 3517.320 2716.890 3518.050 ;
        RECT 2718.010 3517.320 2797.850 3518.050 ;
        RECT 2798.970 3517.320 2878.810 3518.050 ;
        RECT 2879.930 3517.320 2917.220 3518.050 ;
        RECT 2.860 2.680 2917.220 3517.320 ;
        RECT 3.550 1.370 7.950 2.680 ;
        RECT 9.070 1.370 13.930 2.680 ;
        RECT 15.050 1.370 19.910 2.680 ;
        RECT 21.030 1.370 25.890 2.680 ;
        RECT 27.010 1.370 31.870 2.680 ;
        RECT 32.990 1.370 37.850 2.680 ;
        RECT 38.970 1.370 43.370 2.680 ;
        RECT 44.490 1.370 49.350 2.680 ;
        RECT 50.470 1.370 55.330 2.680 ;
        RECT 56.450 1.370 61.310 2.680 ;
        RECT 62.430 1.370 67.290 2.680 ;
        RECT 68.410 1.370 73.270 2.680 ;
        RECT 74.390 1.370 79.250 2.680 ;
        RECT 80.370 1.370 84.770 2.680 ;
        RECT 85.890 1.370 90.750 2.680 ;
        RECT 91.870 1.370 96.730 2.680 ;
        RECT 97.850 1.370 102.710 2.680 ;
        RECT 103.830 1.370 108.690 2.680 ;
        RECT 109.810 1.370 114.670 2.680 ;
        RECT 115.790 1.370 120.650 2.680 ;
        RECT 121.770 1.370 126.170 2.680 ;
        RECT 127.290 1.370 132.150 2.680 ;
        RECT 133.270 1.370 138.130 2.680 ;
        RECT 139.250 1.370 144.110 2.680 ;
        RECT 145.230 1.370 150.090 2.680 ;
        RECT 151.210 1.370 156.070 2.680 ;
        RECT 157.190 1.370 161.590 2.680 ;
        RECT 162.710 1.370 167.570 2.680 ;
        RECT 168.690 1.370 173.550 2.680 ;
        RECT 174.670 1.370 179.530 2.680 ;
        RECT 180.650 1.370 185.510 2.680 ;
        RECT 186.630 1.370 191.490 2.680 ;
        RECT 192.610 1.370 197.470 2.680 ;
        RECT 198.590 1.370 202.990 2.680 ;
        RECT 204.110 1.370 208.970 2.680 ;
        RECT 210.090 1.370 214.950 2.680 ;
        RECT 216.070 1.370 220.930 2.680 ;
        RECT 222.050 1.370 226.910 2.680 ;
        RECT 228.030 1.370 232.890 2.680 ;
        RECT 234.010 1.370 238.870 2.680 ;
        RECT 239.990 1.370 244.390 2.680 ;
        RECT 245.510 1.370 250.370 2.680 ;
        RECT 251.490 1.370 256.350 2.680 ;
        RECT 257.470 1.370 262.330 2.680 ;
        RECT 263.450 1.370 268.310 2.680 ;
        RECT 269.430 1.370 274.290 2.680 ;
        RECT 275.410 1.370 279.810 2.680 ;
        RECT 280.930 1.370 285.790 2.680 ;
        RECT 286.910 1.370 291.770 2.680 ;
        RECT 292.890 1.370 297.750 2.680 ;
        RECT 298.870 1.370 303.730 2.680 ;
        RECT 304.850 1.370 309.710 2.680 ;
        RECT 310.830 1.370 315.690 2.680 ;
        RECT 316.810 1.370 321.210 2.680 ;
        RECT 322.330 1.370 327.190 2.680 ;
        RECT 328.310 1.370 333.170 2.680 ;
        RECT 334.290 1.370 339.150 2.680 ;
        RECT 340.270 1.370 345.130 2.680 ;
        RECT 346.250 1.370 351.110 2.680 ;
        RECT 352.230 1.370 357.090 2.680 ;
        RECT 358.210 1.370 362.610 2.680 ;
        RECT 363.730 1.370 368.590 2.680 ;
        RECT 369.710 1.370 374.570 2.680 ;
        RECT 375.690 1.370 380.550 2.680 ;
        RECT 381.670 1.370 386.530 2.680 ;
        RECT 387.650 1.370 392.510 2.680 ;
        RECT 393.630 1.370 398.030 2.680 ;
        RECT 399.150 1.370 404.010 2.680 ;
        RECT 405.130 1.370 409.990 2.680 ;
        RECT 411.110 1.370 415.970 2.680 ;
        RECT 417.090 1.370 421.950 2.680 ;
        RECT 423.070 1.370 427.930 2.680 ;
        RECT 429.050 1.370 433.910 2.680 ;
        RECT 435.030 1.370 439.430 2.680 ;
        RECT 440.550 1.370 445.410 2.680 ;
        RECT 446.530 1.370 451.390 2.680 ;
        RECT 452.510 1.370 457.370 2.680 ;
        RECT 458.490 1.370 463.350 2.680 ;
        RECT 464.470 1.370 469.330 2.680 ;
        RECT 470.450 1.370 475.310 2.680 ;
        RECT 476.430 1.370 480.830 2.680 ;
        RECT 481.950 1.370 486.810 2.680 ;
        RECT 487.930 1.370 492.790 2.680 ;
        RECT 493.910 1.370 498.770 2.680 ;
        RECT 499.890 1.370 504.750 2.680 ;
        RECT 505.870 1.370 510.730 2.680 ;
        RECT 511.850 1.370 516.250 2.680 ;
        RECT 517.370 1.370 522.230 2.680 ;
        RECT 523.350 1.370 528.210 2.680 ;
        RECT 529.330 1.370 534.190 2.680 ;
        RECT 535.310 1.370 540.170 2.680 ;
        RECT 541.290 1.370 546.150 2.680 ;
        RECT 547.270 1.370 552.130 2.680 ;
        RECT 553.250 1.370 557.650 2.680 ;
        RECT 558.770 1.370 563.630 2.680 ;
        RECT 564.750 1.370 569.610 2.680 ;
        RECT 570.730 1.370 575.590 2.680 ;
        RECT 576.710 1.370 581.570 2.680 ;
        RECT 582.690 1.370 587.550 2.680 ;
        RECT 588.670 1.370 593.530 2.680 ;
        RECT 594.650 1.370 599.050 2.680 ;
        RECT 600.170 1.370 605.030 2.680 ;
        RECT 606.150 1.370 611.010 2.680 ;
        RECT 612.130 1.370 616.990 2.680 ;
        RECT 618.110 1.370 622.970 2.680 ;
        RECT 624.090 1.370 628.950 2.680 ;
        RECT 630.070 1.370 634.470 2.680 ;
        RECT 635.590 1.370 640.450 2.680 ;
        RECT 641.570 1.370 646.430 2.680 ;
        RECT 647.550 1.370 652.410 2.680 ;
        RECT 653.530 1.370 658.390 2.680 ;
        RECT 659.510 1.370 664.370 2.680 ;
        RECT 665.490 1.370 670.350 2.680 ;
        RECT 671.470 1.370 675.870 2.680 ;
        RECT 676.990 1.370 681.850 2.680 ;
        RECT 682.970 1.370 687.830 2.680 ;
        RECT 688.950 1.370 693.810 2.680 ;
        RECT 694.930 1.370 699.790 2.680 ;
        RECT 700.910 1.370 705.770 2.680 ;
        RECT 706.890 1.370 711.750 2.680 ;
        RECT 712.870 1.370 717.270 2.680 ;
        RECT 718.390 1.370 723.250 2.680 ;
        RECT 724.370 1.370 729.230 2.680 ;
        RECT 730.350 1.370 735.210 2.680 ;
        RECT 736.330 1.370 741.190 2.680 ;
        RECT 742.310 1.370 747.170 2.680 ;
        RECT 748.290 1.370 752.690 2.680 ;
        RECT 753.810 1.370 758.670 2.680 ;
        RECT 759.790 1.370 764.650 2.680 ;
        RECT 765.770 1.370 770.630 2.680 ;
        RECT 771.750 1.370 776.610 2.680 ;
        RECT 777.730 1.370 782.590 2.680 ;
        RECT 783.710 1.370 788.570 2.680 ;
        RECT 789.690 1.370 794.090 2.680 ;
        RECT 795.210 1.370 800.070 2.680 ;
        RECT 801.190 1.370 806.050 2.680 ;
        RECT 807.170 1.370 812.030 2.680 ;
        RECT 813.150 1.370 818.010 2.680 ;
        RECT 819.130 1.370 823.990 2.680 ;
        RECT 825.110 1.370 829.970 2.680 ;
        RECT 831.090 1.370 835.490 2.680 ;
        RECT 836.610 1.370 841.470 2.680 ;
        RECT 842.590 1.370 847.450 2.680 ;
        RECT 848.570 1.370 853.430 2.680 ;
        RECT 854.550 1.370 859.410 2.680 ;
        RECT 860.530 1.370 865.390 2.680 ;
        RECT 866.510 1.370 870.910 2.680 ;
        RECT 872.030 1.370 876.890 2.680 ;
        RECT 878.010 1.370 882.870 2.680 ;
        RECT 883.990 1.370 888.850 2.680 ;
        RECT 889.970 1.370 894.830 2.680 ;
        RECT 895.950 1.370 900.810 2.680 ;
        RECT 901.930 1.370 906.790 2.680 ;
        RECT 907.910 1.370 912.310 2.680 ;
        RECT 913.430 1.370 918.290 2.680 ;
        RECT 919.410 1.370 924.270 2.680 ;
        RECT 925.390 1.370 930.250 2.680 ;
        RECT 931.370 1.370 936.230 2.680 ;
        RECT 937.350 1.370 942.210 2.680 ;
        RECT 943.330 1.370 948.190 2.680 ;
        RECT 949.310 1.370 953.710 2.680 ;
        RECT 954.830 1.370 959.690 2.680 ;
        RECT 960.810 1.370 965.670 2.680 ;
        RECT 966.790 1.370 971.650 2.680 ;
        RECT 972.770 1.370 977.630 2.680 ;
        RECT 978.750 1.370 983.610 2.680 ;
        RECT 984.730 1.370 989.130 2.680 ;
        RECT 990.250 1.370 995.110 2.680 ;
        RECT 996.230 1.370 1001.090 2.680 ;
        RECT 1002.210 1.370 1007.070 2.680 ;
        RECT 1008.190 1.370 1013.050 2.680 ;
        RECT 1014.170 1.370 1019.030 2.680 ;
        RECT 1020.150 1.370 1025.010 2.680 ;
        RECT 1026.130 1.370 1030.530 2.680 ;
        RECT 1031.650 1.370 1036.510 2.680 ;
        RECT 1037.630 1.370 1042.490 2.680 ;
        RECT 1043.610 1.370 1048.470 2.680 ;
        RECT 1049.590 1.370 1054.450 2.680 ;
        RECT 1055.570 1.370 1060.430 2.680 ;
        RECT 1061.550 1.370 1066.410 2.680 ;
        RECT 1067.530 1.370 1071.930 2.680 ;
        RECT 1073.050 1.370 1077.910 2.680 ;
        RECT 1079.030 1.370 1083.890 2.680 ;
        RECT 1085.010 1.370 1089.870 2.680 ;
        RECT 1090.990 1.370 1095.850 2.680 ;
        RECT 1096.970 1.370 1101.830 2.680 ;
        RECT 1102.950 1.370 1107.350 2.680 ;
        RECT 1108.470 1.370 1113.330 2.680 ;
        RECT 1114.450 1.370 1119.310 2.680 ;
        RECT 1120.430 1.370 1125.290 2.680 ;
        RECT 1126.410 1.370 1131.270 2.680 ;
        RECT 1132.390 1.370 1137.250 2.680 ;
        RECT 1138.370 1.370 1143.230 2.680 ;
        RECT 1144.350 1.370 1148.750 2.680 ;
        RECT 1149.870 1.370 1154.730 2.680 ;
        RECT 1155.850 1.370 1160.710 2.680 ;
        RECT 1161.830 1.370 1166.690 2.680 ;
        RECT 1167.810 1.370 1172.670 2.680 ;
        RECT 1173.790 1.370 1178.650 2.680 ;
        RECT 1179.770 1.370 1184.630 2.680 ;
        RECT 1185.750 1.370 1190.150 2.680 ;
        RECT 1191.270 1.370 1196.130 2.680 ;
        RECT 1197.250 1.370 1202.110 2.680 ;
        RECT 1203.230 1.370 1208.090 2.680 ;
        RECT 1209.210 1.370 1214.070 2.680 ;
        RECT 1215.190 1.370 1220.050 2.680 ;
        RECT 1221.170 1.370 1225.570 2.680 ;
        RECT 1226.690 1.370 1231.550 2.680 ;
        RECT 1232.670 1.370 1237.530 2.680 ;
        RECT 1238.650 1.370 1243.510 2.680 ;
        RECT 1244.630 1.370 1249.490 2.680 ;
        RECT 1250.610 1.370 1255.470 2.680 ;
        RECT 1256.590 1.370 1261.450 2.680 ;
        RECT 1262.570 1.370 1266.970 2.680 ;
        RECT 1268.090 1.370 1272.950 2.680 ;
        RECT 1274.070 1.370 1278.930 2.680 ;
        RECT 1280.050 1.370 1284.910 2.680 ;
        RECT 1286.030 1.370 1290.890 2.680 ;
        RECT 1292.010 1.370 1296.870 2.680 ;
        RECT 1297.990 1.370 1302.850 2.680 ;
        RECT 1303.970 1.370 1308.370 2.680 ;
        RECT 1309.490 1.370 1314.350 2.680 ;
        RECT 1315.470 1.370 1320.330 2.680 ;
        RECT 1321.450 1.370 1326.310 2.680 ;
        RECT 1327.430 1.370 1332.290 2.680 ;
        RECT 1333.410 1.370 1338.270 2.680 ;
        RECT 1339.390 1.370 1343.790 2.680 ;
        RECT 1344.910 1.370 1349.770 2.680 ;
        RECT 1350.890 1.370 1355.750 2.680 ;
        RECT 1356.870 1.370 1361.730 2.680 ;
        RECT 1362.850 1.370 1367.710 2.680 ;
        RECT 1368.830 1.370 1373.690 2.680 ;
        RECT 1374.810 1.370 1379.670 2.680 ;
        RECT 1380.790 1.370 1385.190 2.680 ;
        RECT 1386.310 1.370 1391.170 2.680 ;
        RECT 1392.290 1.370 1397.150 2.680 ;
        RECT 1398.270 1.370 1403.130 2.680 ;
        RECT 1404.250 1.370 1409.110 2.680 ;
        RECT 1410.230 1.370 1415.090 2.680 ;
        RECT 1416.210 1.370 1421.070 2.680 ;
        RECT 1422.190 1.370 1426.590 2.680 ;
        RECT 1427.710 1.370 1432.570 2.680 ;
        RECT 1433.690 1.370 1438.550 2.680 ;
        RECT 1439.670 1.370 1444.530 2.680 ;
        RECT 1445.650 1.370 1450.510 2.680 ;
        RECT 1451.630 1.370 1456.490 2.680 ;
        RECT 1457.610 1.370 1462.470 2.680 ;
        RECT 1463.590 1.370 1467.990 2.680 ;
        RECT 1469.110 1.370 1473.970 2.680 ;
        RECT 1475.090 1.370 1479.950 2.680 ;
        RECT 1481.070 1.370 1485.930 2.680 ;
        RECT 1487.050 1.370 1491.910 2.680 ;
        RECT 1493.030 1.370 1497.890 2.680 ;
        RECT 1499.010 1.370 1503.410 2.680 ;
        RECT 1504.530 1.370 1509.390 2.680 ;
        RECT 1510.510 1.370 1515.370 2.680 ;
        RECT 1516.490 1.370 1521.350 2.680 ;
        RECT 1522.470 1.370 1527.330 2.680 ;
        RECT 1528.450 1.370 1533.310 2.680 ;
        RECT 1534.430 1.370 1539.290 2.680 ;
        RECT 1540.410 1.370 1544.810 2.680 ;
        RECT 1545.930 1.370 1550.790 2.680 ;
        RECT 1551.910 1.370 1556.770 2.680 ;
        RECT 1557.890 1.370 1562.750 2.680 ;
        RECT 1563.870 1.370 1568.730 2.680 ;
        RECT 1569.850 1.370 1574.710 2.680 ;
        RECT 1575.830 1.370 1580.690 2.680 ;
        RECT 1581.810 1.370 1586.210 2.680 ;
        RECT 1587.330 1.370 1592.190 2.680 ;
        RECT 1593.310 1.370 1598.170 2.680 ;
        RECT 1599.290 1.370 1604.150 2.680 ;
        RECT 1605.270 1.370 1610.130 2.680 ;
        RECT 1611.250 1.370 1616.110 2.680 ;
        RECT 1617.230 1.370 1621.630 2.680 ;
        RECT 1622.750 1.370 1627.610 2.680 ;
        RECT 1628.730 1.370 1633.590 2.680 ;
        RECT 1634.710 1.370 1639.570 2.680 ;
        RECT 1640.690 1.370 1645.550 2.680 ;
        RECT 1646.670 1.370 1651.530 2.680 ;
        RECT 1652.650 1.370 1657.510 2.680 ;
        RECT 1658.630 1.370 1663.030 2.680 ;
        RECT 1664.150 1.370 1669.010 2.680 ;
        RECT 1670.130 1.370 1674.990 2.680 ;
        RECT 1676.110 1.370 1680.970 2.680 ;
        RECT 1682.090 1.370 1686.950 2.680 ;
        RECT 1688.070 1.370 1692.930 2.680 ;
        RECT 1694.050 1.370 1698.910 2.680 ;
        RECT 1700.030 1.370 1704.430 2.680 ;
        RECT 1705.550 1.370 1710.410 2.680 ;
        RECT 1711.530 1.370 1716.390 2.680 ;
        RECT 1717.510 1.370 1722.370 2.680 ;
        RECT 1723.490 1.370 1728.350 2.680 ;
        RECT 1729.470 1.370 1734.330 2.680 ;
        RECT 1735.450 1.370 1739.850 2.680 ;
        RECT 1740.970 1.370 1745.830 2.680 ;
        RECT 1746.950 1.370 1751.810 2.680 ;
        RECT 1752.930 1.370 1757.790 2.680 ;
        RECT 1758.910 1.370 1763.770 2.680 ;
        RECT 1764.890 1.370 1769.750 2.680 ;
        RECT 1770.870 1.370 1775.730 2.680 ;
        RECT 1776.850 1.370 1781.250 2.680 ;
        RECT 1782.370 1.370 1787.230 2.680 ;
        RECT 1788.350 1.370 1793.210 2.680 ;
        RECT 1794.330 1.370 1799.190 2.680 ;
        RECT 1800.310 1.370 1805.170 2.680 ;
        RECT 1806.290 1.370 1811.150 2.680 ;
        RECT 1812.270 1.370 1817.130 2.680 ;
        RECT 1818.250 1.370 1822.650 2.680 ;
        RECT 1823.770 1.370 1828.630 2.680 ;
        RECT 1829.750 1.370 1834.610 2.680 ;
        RECT 1835.730 1.370 1840.590 2.680 ;
        RECT 1841.710 1.370 1846.570 2.680 ;
        RECT 1847.690 1.370 1852.550 2.680 ;
        RECT 1853.670 1.370 1858.070 2.680 ;
        RECT 1859.190 1.370 1864.050 2.680 ;
        RECT 1865.170 1.370 1870.030 2.680 ;
        RECT 1871.150 1.370 1876.010 2.680 ;
        RECT 1877.130 1.370 1881.990 2.680 ;
        RECT 1883.110 1.370 1887.970 2.680 ;
        RECT 1889.090 1.370 1893.950 2.680 ;
        RECT 1895.070 1.370 1899.470 2.680 ;
        RECT 1900.590 1.370 1905.450 2.680 ;
        RECT 1906.570 1.370 1911.430 2.680 ;
        RECT 1912.550 1.370 1917.410 2.680 ;
        RECT 1918.530 1.370 1923.390 2.680 ;
        RECT 1924.510 1.370 1929.370 2.680 ;
        RECT 1930.490 1.370 1935.350 2.680 ;
        RECT 1936.470 1.370 1940.870 2.680 ;
        RECT 1941.990 1.370 1946.850 2.680 ;
        RECT 1947.970 1.370 1952.830 2.680 ;
        RECT 1953.950 1.370 1958.810 2.680 ;
        RECT 1959.930 1.370 1964.790 2.680 ;
        RECT 1965.910 1.370 1970.770 2.680 ;
        RECT 1971.890 1.370 1976.290 2.680 ;
        RECT 1977.410 1.370 1982.270 2.680 ;
        RECT 1983.390 1.370 1988.250 2.680 ;
        RECT 1989.370 1.370 1994.230 2.680 ;
        RECT 1995.350 1.370 2000.210 2.680 ;
        RECT 2001.330 1.370 2006.190 2.680 ;
        RECT 2007.310 1.370 2012.170 2.680 ;
        RECT 2013.290 1.370 2017.690 2.680 ;
        RECT 2018.810 1.370 2023.670 2.680 ;
        RECT 2024.790 1.370 2029.650 2.680 ;
        RECT 2030.770 1.370 2035.630 2.680 ;
        RECT 2036.750 1.370 2041.610 2.680 ;
        RECT 2042.730 1.370 2047.590 2.680 ;
        RECT 2048.710 1.370 2053.570 2.680 ;
        RECT 2054.690 1.370 2059.090 2.680 ;
        RECT 2060.210 1.370 2065.070 2.680 ;
        RECT 2066.190 1.370 2071.050 2.680 ;
        RECT 2072.170 1.370 2077.030 2.680 ;
        RECT 2078.150 1.370 2083.010 2.680 ;
        RECT 2084.130 1.370 2088.990 2.680 ;
        RECT 2090.110 1.370 2094.510 2.680 ;
        RECT 2095.630 1.370 2100.490 2.680 ;
        RECT 2101.610 1.370 2106.470 2.680 ;
        RECT 2107.590 1.370 2112.450 2.680 ;
        RECT 2113.570 1.370 2118.430 2.680 ;
        RECT 2119.550 1.370 2124.410 2.680 ;
        RECT 2125.530 1.370 2130.390 2.680 ;
        RECT 2131.510 1.370 2135.910 2.680 ;
        RECT 2137.030 1.370 2141.890 2.680 ;
        RECT 2143.010 1.370 2147.870 2.680 ;
        RECT 2148.990 1.370 2153.850 2.680 ;
        RECT 2154.970 1.370 2159.830 2.680 ;
        RECT 2160.950 1.370 2165.810 2.680 ;
        RECT 2166.930 1.370 2171.790 2.680 ;
        RECT 2172.910 1.370 2177.310 2.680 ;
        RECT 2178.430 1.370 2183.290 2.680 ;
        RECT 2184.410 1.370 2189.270 2.680 ;
        RECT 2190.390 1.370 2195.250 2.680 ;
        RECT 2196.370 1.370 2201.230 2.680 ;
        RECT 2202.350 1.370 2207.210 2.680 ;
        RECT 2208.330 1.370 2212.730 2.680 ;
        RECT 2213.850 1.370 2218.710 2.680 ;
        RECT 2219.830 1.370 2224.690 2.680 ;
        RECT 2225.810 1.370 2230.670 2.680 ;
        RECT 2231.790 1.370 2236.650 2.680 ;
        RECT 2237.770 1.370 2242.630 2.680 ;
        RECT 2243.750 1.370 2248.610 2.680 ;
        RECT 2249.730 1.370 2254.130 2.680 ;
        RECT 2255.250 1.370 2260.110 2.680 ;
        RECT 2261.230 1.370 2266.090 2.680 ;
        RECT 2267.210 1.370 2272.070 2.680 ;
        RECT 2273.190 1.370 2278.050 2.680 ;
        RECT 2279.170 1.370 2284.030 2.680 ;
        RECT 2285.150 1.370 2290.010 2.680 ;
        RECT 2291.130 1.370 2295.530 2.680 ;
        RECT 2296.650 1.370 2301.510 2.680 ;
        RECT 2302.630 1.370 2307.490 2.680 ;
        RECT 2308.610 1.370 2313.470 2.680 ;
        RECT 2314.590 1.370 2319.450 2.680 ;
        RECT 2320.570 1.370 2325.430 2.680 ;
        RECT 2326.550 1.370 2330.950 2.680 ;
        RECT 2332.070 1.370 2336.930 2.680 ;
        RECT 2338.050 1.370 2342.910 2.680 ;
        RECT 2344.030 1.370 2348.890 2.680 ;
        RECT 2350.010 1.370 2354.870 2.680 ;
        RECT 2355.990 1.370 2360.850 2.680 ;
        RECT 2361.970 1.370 2366.830 2.680 ;
        RECT 2367.950 1.370 2372.350 2.680 ;
        RECT 2373.470 1.370 2378.330 2.680 ;
        RECT 2379.450 1.370 2384.310 2.680 ;
        RECT 2385.430 1.370 2390.290 2.680 ;
        RECT 2391.410 1.370 2396.270 2.680 ;
        RECT 2397.390 1.370 2402.250 2.680 ;
        RECT 2403.370 1.370 2408.230 2.680 ;
        RECT 2409.350 1.370 2413.750 2.680 ;
        RECT 2414.870 1.370 2419.730 2.680 ;
        RECT 2420.850 1.370 2425.710 2.680 ;
        RECT 2426.830 1.370 2431.690 2.680 ;
        RECT 2432.810 1.370 2437.670 2.680 ;
        RECT 2438.790 1.370 2443.650 2.680 ;
        RECT 2444.770 1.370 2449.170 2.680 ;
        RECT 2450.290 1.370 2455.150 2.680 ;
        RECT 2456.270 1.370 2461.130 2.680 ;
        RECT 2462.250 1.370 2467.110 2.680 ;
        RECT 2468.230 1.370 2473.090 2.680 ;
        RECT 2474.210 1.370 2479.070 2.680 ;
        RECT 2480.190 1.370 2485.050 2.680 ;
        RECT 2486.170 1.370 2490.570 2.680 ;
        RECT 2491.690 1.370 2496.550 2.680 ;
        RECT 2497.670 1.370 2502.530 2.680 ;
        RECT 2503.650 1.370 2508.510 2.680 ;
        RECT 2509.630 1.370 2514.490 2.680 ;
        RECT 2515.610 1.370 2520.470 2.680 ;
        RECT 2521.590 1.370 2526.450 2.680 ;
        RECT 2527.570 1.370 2531.970 2.680 ;
        RECT 2533.090 1.370 2537.950 2.680 ;
        RECT 2539.070 1.370 2543.930 2.680 ;
        RECT 2545.050 1.370 2549.910 2.680 ;
        RECT 2551.030 1.370 2555.890 2.680 ;
        RECT 2557.010 1.370 2561.870 2.680 ;
        RECT 2562.990 1.370 2567.390 2.680 ;
        RECT 2568.510 1.370 2573.370 2.680 ;
        RECT 2574.490 1.370 2579.350 2.680 ;
        RECT 2580.470 1.370 2585.330 2.680 ;
        RECT 2586.450 1.370 2591.310 2.680 ;
        RECT 2592.430 1.370 2597.290 2.680 ;
        RECT 2598.410 1.370 2603.270 2.680 ;
        RECT 2604.390 1.370 2608.790 2.680 ;
        RECT 2609.910 1.370 2614.770 2.680 ;
        RECT 2615.890 1.370 2620.750 2.680 ;
        RECT 2621.870 1.370 2626.730 2.680 ;
        RECT 2627.850 1.370 2632.710 2.680 ;
        RECT 2633.830 1.370 2638.690 2.680 ;
        RECT 2639.810 1.370 2644.670 2.680 ;
        RECT 2645.790 1.370 2650.190 2.680 ;
        RECT 2651.310 1.370 2656.170 2.680 ;
        RECT 2657.290 1.370 2662.150 2.680 ;
        RECT 2663.270 1.370 2668.130 2.680 ;
        RECT 2669.250 1.370 2674.110 2.680 ;
        RECT 2675.230 1.370 2680.090 2.680 ;
        RECT 2681.210 1.370 2685.610 2.680 ;
        RECT 2686.730 1.370 2691.590 2.680 ;
        RECT 2692.710 1.370 2697.570 2.680 ;
        RECT 2698.690 1.370 2703.550 2.680 ;
        RECT 2704.670 1.370 2709.530 2.680 ;
        RECT 2710.650 1.370 2715.510 2.680 ;
        RECT 2716.630 1.370 2721.490 2.680 ;
        RECT 2722.610 1.370 2727.010 2.680 ;
        RECT 2728.130 1.370 2732.990 2.680 ;
        RECT 2734.110 1.370 2738.970 2.680 ;
        RECT 2740.090 1.370 2744.950 2.680 ;
        RECT 2746.070 1.370 2750.930 2.680 ;
        RECT 2752.050 1.370 2756.910 2.680 ;
        RECT 2758.030 1.370 2762.890 2.680 ;
        RECT 2764.010 1.370 2768.410 2.680 ;
        RECT 2769.530 1.370 2774.390 2.680 ;
        RECT 2775.510 1.370 2780.370 2.680 ;
        RECT 2781.490 1.370 2786.350 2.680 ;
        RECT 2787.470 1.370 2792.330 2.680 ;
        RECT 2793.450 1.370 2798.310 2.680 ;
        RECT 2799.430 1.370 2803.830 2.680 ;
        RECT 2804.950 1.370 2809.810 2.680 ;
        RECT 2810.930 1.370 2815.790 2.680 ;
        RECT 2816.910 1.370 2821.770 2.680 ;
        RECT 2822.890 1.370 2827.750 2.680 ;
        RECT 2828.870 1.370 2833.730 2.680 ;
        RECT 2834.850 1.370 2839.710 2.680 ;
        RECT 2840.830 1.370 2845.230 2.680 ;
        RECT 2846.350 1.370 2851.210 2.680 ;
        RECT 2852.330 1.370 2857.190 2.680 ;
        RECT 2858.310 1.370 2863.170 2.680 ;
        RECT 2864.290 1.370 2869.150 2.680 ;
        RECT 2870.270 1.370 2875.130 2.680 ;
        RECT 2876.250 1.370 2881.110 2.680 ;
        RECT 2882.230 1.370 2886.630 2.680 ;
        RECT 2887.750 1.370 2892.610 2.680 ;
        RECT 2893.730 1.370 2898.590 2.680 ;
        RECT 2899.710 1.370 2904.570 2.680 ;
        RECT 2905.690 1.370 2910.550 2.680 ;
        RECT 2911.670 1.370 2916.530 2.680 ;
      LAYER met3 ;
        RECT 2.400 3487.700 2917.600 3508.965 ;
        RECT 2.800 3487.020 2917.600 3487.700 ;
        RECT 2.800 3485.700 2917.200 3487.020 ;
        RECT 2.400 3485.020 2917.200 3485.700 ;
        RECT 2.400 3422.420 2917.600 3485.020 ;
        RECT 2.800 3420.420 2917.600 3422.420 ;
        RECT 2.400 3420.380 2917.600 3420.420 ;
        RECT 2.400 3418.380 2917.200 3420.380 ;
        RECT 2.400 3357.140 2917.600 3418.380 ;
        RECT 2.800 3355.140 2917.600 3357.140 ;
        RECT 2.400 3354.420 2917.600 3355.140 ;
        RECT 2.400 3352.420 2917.200 3354.420 ;
        RECT 2.400 3291.860 2917.600 3352.420 ;
        RECT 2.800 3289.860 2917.600 3291.860 ;
        RECT 2.400 3287.780 2917.600 3289.860 ;
        RECT 2.400 3285.780 2917.200 3287.780 ;
        RECT 2.400 3226.580 2917.600 3285.780 ;
        RECT 2.800 3224.580 2917.600 3226.580 ;
        RECT 2.400 3221.140 2917.600 3224.580 ;
        RECT 2.400 3219.140 2917.200 3221.140 ;
        RECT 2.400 3161.300 2917.600 3219.140 ;
        RECT 2.800 3159.300 2917.600 3161.300 ;
        RECT 2.400 3155.180 2917.600 3159.300 ;
        RECT 2.400 3153.180 2917.200 3155.180 ;
        RECT 2.400 3096.700 2917.600 3153.180 ;
        RECT 2.800 3094.700 2917.600 3096.700 ;
        RECT 2.400 3088.540 2917.600 3094.700 ;
        RECT 2.400 3086.540 2917.200 3088.540 ;
        RECT 2.400 3031.420 2917.600 3086.540 ;
        RECT 2.800 3029.420 2917.600 3031.420 ;
        RECT 2.400 3021.900 2917.600 3029.420 ;
        RECT 2.400 3019.900 2917.200 3021.900 ;
        RECT 2.400 2966.140 2917.600 3019.900 ;
        RECT 2.800 2964.140 2917.600 2966.140 ;
        RECT 2.400 2955.940 2917.600 2964.140 ;
        RECT 2.400 2953.940 2917.200 2955.940 ;
        RECT 2.400 2900.860 2917.600 2953.940 ;
        RECT 2.800 2898.860 2917.600 2900.860 ;
        RECT 2.400 2889.300 2917.600 2898.860 ;
        RECT 2.400 2887.300 2917.200 2889.300 ;
        RECT 2.400 2835.580 2917.600 2887.300 ;
        RECT 2.800 2833.580 2917.600 2835.580 ;
        RECT 2.400 2822.660 2917.600 2833.580 ;
        RECT 2.400 2820.660 2917.200 2822.660 ;
        RECT 2.400 2770.300 2917.600 2820.660 ;
        RECT 2.800 2768.300 2917.600 2770.300 ;
        RECT 2.400 2756.700 2917.600 2768.300 ;
        RECT 2.400 2754.700 2917.200 2756.700 ;
        RECT 2.400 2705.020 2917.600 2754.700 ;
        RECT 2.800 2703.020 2917.600 2705.020 ;
        RECT 2.400 2690.060 2917.600 2703.020 ;
        RECT 2.400 2688.060 2917.200 2690.060 ;
        RECT 2.400 2640.420 2917.600 2688.060 ;
        RECT 2.800 2638.420 2917.600 2640.420 ;
        RECT 2.400 2623.420 2917.600 2638.420 ;
        RECT 2.400 2621.420 2917.200 2623.420 ;
        RECT 2.400 2575.140 2917.600 2621.420 ;
        RECT 2.800 2573.140 2917.600 2575.140 ;
        RECT 2.400 2557.460 2917.600 2573.140 ;
        RECT 2.400 2555.460 2917.200 2557.460 ;
        RECT 2.400 2509.860 2917.600 2555.460 ;
        RECT 2.800 2507.860 2917.600 2509.860 ;
        RECT 2.400 2490.820 2917.600 2507.860 ;
        RECT 2.400 2488.820 2917.200 2490.820 ;
        RECT 2.400 2444.580 2917.600 2488.820 ;
        RECT 2.800 2442.580 2917.600 2444.580 ;
        RECT 2.400 2424.180 2917.600 2442.580 ;
        RECT 2.400 2422.180 2917.200 2424.180 ;
        RECT 2.400 2379.300 2917.600 2422.180 ;
        RECT 2.800 2377.300 2917.600 2379.300 ;
        RECT 2.400 2358.220 2917.600 2377.300 ;
        RECT 2.400 2356.220 2917.200 2358.220 ;
        RECT 2.400 2314.020 2917.600 2356.220 ;
        RECT 2.800 2312.020 2917.600 2314.020 ;
        RECT 2.400 2291.580 2917.600 2312.020 ;
        RECT 2.400 2289.580 2917.200 2291.580 ;
        RECT 2.400 2248.740 2917.600 2289.580 ;
        RECT 2.800 2246.740 2917.600 2248.740 ;
        RECT 2.400 2224.940 2917.600 2246.740 ;
        RECT 2.400 2222.940 2917.200 2224.940 ;
        RECT 2.400 2184.140 2917.600 2222.940 ;
        RECT 2.800 2182.140 2917.600 2184.140 ;
        RECT 2.400 2158.980 2917.600 2182.140 ;
        RECT 2.400 2156.980 2917.200 2158.980 ;
        RECT 2.400 2118.860 2917.600 2156.980 ;
        RECT 2.800 2116.860 2917.600 2118.860 ;
        RECT 2.400 2092.340 2917.600 2116.860 ;
        RECT 2.400 2090.340 2917.200 2092.340 ;
        RECT 2.400 2053.580 2917.600 2090.340 ;
        RECT 2.800 2051.580 2917.600 2053.580 ;
        RECT 2.400 2025.700 2917.600 2051.580 ;
        RECT 2.400 2023.700 2917.200 2025.700 ;
        RECT 2.400 1988.300 2917.600 2023.700 ;
        RECT 2.800 1986.300 2917.600 1988.300 ;
        RECT 2.400 1959.740 2917.600 1986.300 ;
        RECT 2.400 1957.740 2917.200 1959.740 ;
        RECT 2.400 1923.020 2917.600 1957.740 ;
        RECT 2.800 1921.020 2917.600 1923.020 ;
        RECT 2.400 1893.100 2917.600 1921.020 ;
        RECT 2.400 1891.100 2917.200 1893.100 ;
        RECT 2.400 1857.740 2917.600 1891.100 ;
        RECT 2.800 1855.740 2917.600 1857.740 ;
        RECT 2.400 1826.460 2917.600 1855.740 ;
        RECT 2.400 1824.460 2917.200 1826.460 ;
        RECT 2.400 1793.140 2917.600 1824.460 ;
        RECT 2.800 1791.140 2917.600 1793.140 ;
        RECT 2.400 1760.500 2917.600 1791.140 ;
        RECT 2.400 1758.500 2917.200 1760.500 ;
        RECT 2.400 1727.860 2917.600 1758.500 ;
        RECT 2.800 1725.860 2917.600 1727.860 ;
        RECT 2.400 1693.860 2917.600 1725.860 ;
        RECT 2.400 1691.860 2917.200 1693.860 ;
        RECT 2.400 1662.580 2917.600 1691.860 ;
        RECT 2.800 1660.580 2917.600 1662.580 ;
        RECT 2.400 1627.220 2917.600 1660.580 ;
        RECT 2.400 1625.220 2917.200 1627.220 ;
        RECT 2.400 1597.300 2917.600 1625.220 ;
        RECT 2.800 1595.300 2917.600 1597.300 ;
        RECT 2.400 1561.260 2917.600 1595.300 ;
        RECT 2.400 1559.260 2917.200 1561.260 ;
        RECT 2.400 1532.020 2917.600 1559.260 ;
        RECT 2.800 1530.020 2917.600 1532.020 ;
        RECT 2.400 1494.620 2917.600 1530.020 ;
        RECT 2.400 1492.620 2917.200 1494.620 ;
        RECT 2.400 1466.740 2917.600 1492.620 ;
        RECT 2.800 1464.740 2917.600 1466.740 ;
        RECT 2.400 1427.980 2917.600 1464.740 ;
        RECT 2.400 1425.980 2917.200 1427.980 ;
        RECT 2.400 1401.460 2917.600 1425.980 ;
        RECT 2.800 1399.460 2917.600 1401.460 ;
        RECT 2.400 1362.020 2917.600 1399.460 ;
        RECT 2.400 1360.020 2917.200 1362.020 ;
        RECT 2.400 1336.860 2917.600 1360.020 ;
        RECT 2.800 1334.860 2917.600 1336.860 ;
        RECT 2.400 1295.380 2917.600 1334.860 ;
        RECT 2.400 1293.380 2917.200 1295.380 ;
        RECT 2.400 1271.580 2917.600 1293.380 ;
        RECT 2.800 1269.580 2917.600 1271.580 ;
        RECT 2.400 1228.740 2917.600 1269.580 ;
        RECT 2.400 1226.740 2917.200 1228.740 ;
        RECT 2.400 1206.300 2917.600 1226.740 ;
        RECT 2.800 1204.300 2917.600 1206.300 ;
        RECT 2.400 1162.780 2917.600 1204.300 ;
        RECT 2.400 1160.780 2917.200 1162.780 ;
        RECT 2.400 1141.020 2917.600 1160.780 ;
        RECT 2.800 1139.020 2917.600 1141.020 ;
        RECT 2.400 1096.140 2917.600 1139.020 ;
        RECT 2.400 1094.140 2917.200 1096.140 ;
        RECT 2.400 1075.740 2917.600 1094.140 ;
        RECT 2.800 1073.740 2917.600 1075.740 ;
        RECT 2.400 1029.500 2917.600 1073.740 ;
        RECT 2.400 1027.500 2917.200 1029.500 ;
        RECT 2.400 1010.460 2917.600 1027.500 ;
        RECT 2.800 1008.460 2917.600 1010.460 ;
        RECT 2.400 963.540 2917.600 1008.460 ;
        RECT 2.400 961.540 2917.200 963.540 ;
        RECT 2.400 945.180 2917.600 961.540 ;
        RECT 2.800 943.180 2917.600 945.180 ;
        RECT 2.400 896.900 2917.600 943.180 ;
        RECT 2.400 894.900 2917.200 896.900 ;
        RECT 2.400 880.580 2917.600 894.900 ;
        RECT 2.800 878.580 2917.600 880.580 ;
        RECT 2.400 830.260 2917.600 878.580 ;
        RECT 2.400 828.260 2917.200 830.260 ;
        RECT 2.400 815.300 2917.600 828.260 ;
        RECT 2.800 813.300 2917.600 815.300 ;
        RECT 2.400 764.300 2917.600 813.300 ;
        RECT 2.400 762.300 2917.200 764.300 ;
        RECT 2.400 750.020 2917.600 762.300 ;
        RECT 2.800 748.020 2917.600 750.020 ;
        RECT 2.400 697.660 2917.600 748.020 ;
        RECT 2.400 695.660 2917.200 697.660 ;
        RECT 2.400 684.740 2917.600 695.660 ;
        RECT 2.800 682.740 2917.600 684.740 ;
        RECT 2.400 631.020 2917.600 682.740 ;
        RECT 2.400 629.020 2917.200 631.020 ;
        RECT 2.400 619.460 2917.600 629.020 ;
        RECT 2.800 617.460 2917.600 619.460 ;
        RECT 2.400 565.060 2917.600 617.460 ;
        RECT 2.400 563.060 2917.200 565.060 ;
        RECT 2.400 554.180 2917.600 563.060 ;
        RECT 2.800 552.180 2917.600 554.180 ;
        RECT 2.400 498.420 2917.600 552.180 ;
        RECT 2.400 496.420 2917.200 498.420 ;
        RECT 2.400 488.900 2917.600 496.420 ;
        RECT 2.800 486.900 2917.600 488.900 ;
        RECT 2.400 431.780 2917.600 486.900 ;
        RECT 2.400 429.780 2917.200 431.780 ;
        RECT 2.400 424.300 2917.600 429.780 ;
        RECT 2.800 422.300 2917.600 424.300 ;
        RECT 2.400 365.820 2917.600 422.300 ;
        RECT 2.400 363.820 2917.200 365.820 ;
        RECT 2.400 359.020 2917.600 363.820 ;
        RECT 2.800 357.020 2917.600 359.020 ;
        RECT 2.400 299.180 2917.600 357.020 ;
        RECT 2.400 297.180 2917.200 299.180 ;
        RECT 2.400 293.740 2917.600 297.180 ;
        RECT 2.800 291.740 2917.600 293.740 ;
        RECT 2.400 232.540 2917.600 291.740 ;
        RECT 2.400 230.540 2917.200 232.540 ;
        RECT 2.400 228.460 2917.600 230.540 ;
        RECT 2.800 226.460 2917.600 228.460 ;
        RECT 2.400 166.580 2917.600 226.460 ;
        RECT 2.400 164.580 2917.200 166.580 ;
        RECT 2.400 163.180 2917.600 164.580 ;
        RECT 2.800 161.180 2917.600 163.180 ;
        RECT 2.400 99.940 2917.600 161.180 ;
        RECT 2.400 97.940 2917.200 99.940 ;
        RECT 2.400 97.900 2917.600 97.940 ;
        RECT 2.800 95.900 2917.600 97.900 ;
        RECT 2.400 33.980 2917.600 95.900 ;
        RECT 2.400 33.300 2917.200 33.980 ;
        RECT 2.800 31.980 2917.200 33.300 ;
        RECT 2.800 31.300 2917.600 31.980 ;
        RECT 2.400 10.715 2917.600 31.300 ;
      LAYER met4 ;
        RECT 178.775 3351.740 188.570 3355.040 ;
        RECT 192.470 3351.980 207.170 3355.040 ;
        RECT 211.070 3351.980 225.770 3355.040 ;
        RECT 229.670 3351.980 244.370 3355.040 ;
        RECT 248.270 3351.980 278.570 3355.040 ;
        RECT 192.470 3351.740 278.570 3351.980 ;
        RECT 282.470 3351.980 297.170 3355.040 ;
        RECT 301.070 3351.980 315.770 3355.040 ;
        RECT 319.670 3351.980 334.370 3355.040 ;
        RECT 338.270 3351.980 368.570 3355.040 ;
        RECT 282.470 3351.740 368.570 3351.980 ;
        RECT 372.470 3351.980 387.170 3355.040 ;
        RECT 391.070 3351.980 405.770 3355.040 ;
        RECT 409.670 3351.980 424.370 3355.040 ;
        RECT 428.270 3351.980 458.570 3355.040 ;
        RECT 372.470 3351.740 458.570 3351.980 ;
        RECT 462.470 3351.980 477.170 3355.040 ;
        RECT 481.070 3351.980 495.770 3355.040 ;
        RECT 499.670 3351.980 514.370 3355.040 ;
        RECT 518.270 3351.980 548.570 3355.040 ;
        RECT 462.470 3351.740 548.570 3351.980 ;
        RECT 552.470 3351.980 567.170 3355.040 ;
        RECT 571.070 3351.980 585.770 3355.040 ;
        RECT 589.670 3351.980 604.370 3355.040 ;
        RECT 608.270 3351.980 638.570 3355.040 ;
        RECT 552.470 3351.740 638.570 3351.980 ;
        RECT 642.470 3351.980 657.170 3355.040 ;
        RECT 661.070 3351.980 675.770 3355.040 ;
        RECT 642.470 3351.740 675.770 3351.980 ;
        RECT 178.775 2885.880 675.770 3351.740 ;
        RECT 178.775 2733.720 188.570 2885.880 ;
        RECT 192.470 2885.640 278.570 2885.880 ;
        RECT 192.470 2733.960 207.170 2885.640 ;
        RECT 211.070 2733.960 225.770 2885.640 ;
        RECT 229.670 2733.960 244.370 2885.640 ;
        RECT 248.270 2733.960 278.570 2885.640 ;
        RECT 192.470 2733.720 278.570 2733.960 ;
        RECT 282.470 2885.640 368.570 2885.880 ;
        RECT 282.470 2733.960 297.170 2885.640 ;
        RECT 301.070 2733.960 315.770 2885.640 ;
        RECT 319.670 2733.960 334.370 2885.640 ;
        RECT 338.270 2733.960 368.570 2885.640 ;
        RECT 282.470 2733.720 368.570 2733.960 ;
        RECT 372.470 2885.640 458.570 2885.880 ;
        RECT 372.470 2733.960 387.170 2885.640 ;
        RECT 391.070 2733.960 405.770 2885.640 ;
        RECT 409.670 2733.960 424.370 2885.640 ;
        RECT 428.270 2733.960 458.570 2885.640 ;
        RECT 372.470 2733.720 458.570 2733.960 ;
        RECT 462.470 2885.640 548.570 2885.880 ;
        RECT 462.470 2733.960 477.170 2885.640 ;
        RECT 481.070 2733.960 495.770 2885.640 ;
        RECT 499.670 2733.960 514.370 2885.640 ;
        RECT 518.270 2733.960 548.570 2885.640 ;
        RECT 462.470 2733.720 548.570 2733.960 ;
        RECT 552.470 2885.640 638.570 2885.880 ;
        RECT 552.470 2733.960 567.170 2885.640 ;
        RECT 571.070 2733.960 585.770 2885.640 ;
        RECT 589.670 2733.960 604.370 2885.640 ;
        RECT 608.270 2733.960 638.570 2885.640 ;
        RECT 552.470 2733.720 638.570 2733.960 ;
        RECT 642.470 2885.640 675.770 2885.880 ;
        RECT 642.470 2733.960 657.170 2885.640 ;
        RECT 661.070 2733.960 675.770 2885.640 ;
        RECT 679.670 2733.960 694.370 3355.040 ;
        RECT 698.270 2733.960 728.570 3355.040 ;
        RECT 642.470 2733.720 728.570 2733.960 ;
        RECT 178.775 2311.380 728.570 2733.720 ;
        RECT 178.775 2156.500 188.570 2311.380 ;
        RECT 192.470 2311.140 278.570 2311.380 ;
        RECT 192.470 2156.740 207.170 2311.140 ;
        RECT 211.070 2156.740 225.770 2311.140 ;
        RECT 229.670 2156.740 244.370 2311.140 ;
        RECT 248.270 2156.740 278.570 2311.140 ;
        RECT 192.470 2156.500 278.570 2156.740 ;
        RECT 282.470 2311.140 368.570 2311.380 ;
        RECT 282.470 2156.740 297.170 2311.140 ;
        RECT 301.070 2156.740 315.770 2311.140 ;
        RECT 319.670 2156.740 334.370 2311.140 ;
        RECT 338.270 2156.740 368.570 2311.140 ;
        RECT 282.470 2156.500 368.570 2156.740 ;
        RECT 372.470 2311.140 458.570 2311.380 ;
        RECT 372.470 2156.740 387.170 2311.140 ;
        RECT 391.070 2156.740 405.770 2311.140 ;
        RECT 409.670 2156.740 424.370 2311.140 ;
        RECT 428.270 2156.740 458.570 2311.140 ;
        RECT 372.470 2156.500 458.570 2156.740 ;
        RECT 462.470 2311.140 548.570 2311.380 ;
        RECT 462.470 2156.740 477.170 2311.140 ;
        RECT 481.070 2156.740 495.770 2311.140 ;
        RECT 499.670 2156.740 514.370 2311.140 ;
        RECT 518.270 2156.740 548.570 2311.140 ;
        RECT 462.470 2156.500 548.570 2156.740 ;
        RECT 552.470 2311.140 638.570 2311.380 ;
        RECT 552.470 2156.740 567.170 2311.140 ;
        RECT 571.070 2156.740 585.770 2311.140 ;
        RECT 589.670 2156.740 604.370 2311.140 ;
        RECT 608.270 2156.740 638.570 2311.140 ;
        RECT 552.470 2156.500 638.570 2156.740 ;
        RECT 642.470 2311.140 728.570 2311.380 ;
        RECT 642.470 2156.740 657.170 2311.140 ;
        RECT 661.070 2156.740 675.770 2311.140 ;
        RECT 679.670 2156.740 694.370 2311.140 ;
        RECT 698.270 2156.740 728.570 2311.140 ;
        RECT 642.470 2156.500 728.570 2156.740 ;
        RECT 732.470 2156.740 747.170 3355.040 ;
        RECT 751.070 2156.740 765.770 3355.040 ;
        RECT 769.670 2156.740 784.370 3355.040 ;
        RECT 788.270 2156.740 818.570 3355.040 ;
        RECT 732.470 2156.500 818.570 2156.740 ;
        RECT 822.470 2156.740 837.170 3355.040 ;
        RECT 841.070 2156.740 855.770 3355.040 ;
        RECT 859.670 2156.740 874.370 3355.040 ;
        RECT 878.270 2156.740 908.570 3355.040 ;
        RECT 822.470 2156.500 908.570 2156.740 ;
        RECT 912.470 2156.500 927.170 3355.040 ;
        RECT 178.775 1465.560 927.170 2156.500 ;
        RECT 178.775 1005.360 188.570 1465.560 ;
        RECT 192.470 1465.320 278.570 1465.560 ;
        RECT 192.470 1005.600 207.170 1465.320 ;
        RECT 211.070 1005.600 225.770 1465.320 ;
        RECT 229.670 1005.600 244.370 1465.320 ;
        RECT 248.270 1005.600 278.570 1465.320 ;
        RECT 192.470 1005.360 278.570 1005.600 ;
        RECT 282.470 1465.320 368.570 1465.560 ;
        RECT 282.470 1005.600 297.170 1465.320 ;
        RECT 301.070 1005.600 315.770 1465.320 ;
        RECT 319.670 1005.600 334.370 1465.320 ;
        RECT 338.270 1005.600 368.570 1465.320 ;
        RECT 282.470 1005.360 368.570 1005.600 ;
        RECT 372.470 1465.320 458.570 1465.560 ;
        RECT 372.470 1005.600 387.170 1465.320 ;
        RECT 391.070 1005.600 405.770 1465.320 ;
        RECT 409.670 1005.600 424.370 1465.320 ;
        RECT 428.270 1005.600 458.570 1465.320 ;
        RECT 372.470 1005.360 458.570 1005.600 ;
        RECT 462.470 1465.320 548.570 1465.560 ;
        RECT 462.470 1005.600 477.170 1465.320 ;
        RECT 481.070 1005.600 495.770 1465.320 ;
        RECT 499.670 1005.600 514.370 1465.320 ;
        RECT 518.270 1005.600 548.570 1465.320 ;
        RECT 462.470 1005.360 548.570 1005.600 ;
        RECT 552.470 1465.320 638.570 1465.560 ;
        RECT 552.470 1005.600 567.170 1465.320 ;
        RECT 571.070 1005.600 585.770 1465.320 ;
        RECT 589.670 1005.600 604.370 1465.320 ;
        RECT 608.270 1005.600 638.570 1465.320 ;
        RECT 552.470 1005.360 638.570 1005.600 ;
        RECT 642.470 1465.320 728.570 1465.560 ;
        RECT 642.470 1005.600 657.170 1465.320 ;
        RECT 661.070 1005.600 675.770 1465.320 ;
        RECT 679.670 1005.600 694.370 1465.320 ;
        RECT 698.270 1005.600 728.570 1465.320 ;
        RECT 642.470 1005.360 728.570 1005.600 ;
        RECT 732.470 1465.320 818.570 1465.560 ;
        RECT 732.470 1005.600 747.170 1465.320 ;
        RECT 751.070 1005.600 765.770 1465.320 ;
        RECT 769.670 1005.600 784.370 1465.320 ;
        RECT 788.270 1005.600 818.570 1465.320 ;
        RECT 732.470 1005.360 818.570 1005.600 ;
        RECT 822.470 1465.320 908.570 1465.560 ;
        RECT 822.470 1005.600 837.170 1465.320 ;
        RECT 841.070 1005.600 855.770 1465.320 ;
        RECT 859.670 1005.600 874.370 1465.320 ;
        RECT 878.270 1005.600 908.570 1465.320 ;
        RECT 822.470 1005.360 908.570 1005.600 ;
        RECT 178.775 568.060 908.570 1005.360 ;
        RECT 178.775 409.780 188.570 568.060 ;
        RECT 192.470 567.820 278.570 568.060 ;
        RECT 192.470 410.020 207.170 567.820 ;
        RECT 211.070 410.020 225.770 567.820 ;
        RECT 229.670 410.020 244.370 567.820 ;
        RECT 248.270 410.020 278.570 567.820 ;
        RECT 192.470 409.780 278.570 410.020 ;
        RECT 282.470 567.820 368.570 568.060 ;
        RECT 282.470 410.020 297.170 567.820 ;
        RECT 301.070 410.020 315.770 567.820 ;
        RECT 319.670 410.020 334.370 567.820 ;
        RECT 338.270 410.020 368.570 567.820 ;
        RECT 282.470 409.780 368.570 410.020 ;
        RECT 372.470 567.820 458.570 568.060 ;
        RECT 372.470 410.020 387.170 567.820 ;
        RECT 391.070 410.020 405.770 567.820 ;
        RECT 409.670 410.020 424.370 567.820 ;
        RECT 428.270 410.020 458.570 567.820 ;
        RECT 372.470 409.780 458.570 410.020 ;
        RECT 462.470 567.820 548.570 568.060 ;
        RECT 462.470 410.020 477.170 567.820 ;
        RECT 481.070 410.020 495.770 567.820 ;
        RECT 499.670 410.020 514.370 567.820 ;
        RECT 518.270 410.020 548.570 567.820 ;
        RECT 462.470 409.780 548.570 410.020 ;
        RECT 552.470 567.820 638.570 568.060 ;
        RECT 552.470 410.020 567.170 567.820 ;
        RECT 571.070 410.020 585.770 567.820 ;
        RECT 589.670 410.020 604.370 567.820 ;
        RECT 608.270 410.020 638.570 567.820 ;
        RECT 552.470 409.780 638.570 410.020 ;
        RECT 642.470 567.820 728.570 568.060 ;
        RECT 642.470 410.020 657.170 567.820 ;
        RECT 661.070 410.020 675.770 567.820 ;
        RECT 679.670 410.020 694.370 567.820 ;
        RECT 642.470 409.780 694.370 410.020 ;
        RECT 178.775 167.640 694.370 409.780 ;
        RECT 178.775 42.335 188.570 167.640 ;
        RECT 192.470 167.400 278.570 167.640 ;
        RECT 192.470 42.335 207.170 167.400 ;
        RECT 211.070 42.335 225.770 167.400 ;
        RECT 229.670 42.335 244.370 167.400 ;
        RECT 248.270 42.335 278.570 167.400 ;
        RECT 282.470 167.400 368.570 167.640 ;
        RECT 282.470 42.335 297.170 167.400 ;
        RECT 301.070 42.335 315.770 167.400 ;
        RECT 319.670 42.335 334.370 167.400 ;
        RECT 338.270 42.335 368.570 167.400 ;
        RECT 372.470 167.400 458.570 167.640 ;
        RECT 372.470 42.335 387.170 167.400 ;
        RECT 391.070 42.335 405.770 167.400 ;
        RECT 409.670 42.335 424.370 167.400 ;
        RECT 428.270 42.335 458.570 167.400 ;
        RECT 462.470 167.400 548.570 167.640 ;
        RECT 462.470 42.335 477.170 167.400 ;
        RECT 481.070 42.335 495.770 167.400 ;
        RECT 499.670 42.335 514.370 167.400 ;
        RECT 518.270 42.335 548.570 167.400 ;
        RECT 552.470 167.400 638.570 167.640 ;
        RECT 552.470 42.335 567.170 167.400 ;
        RECT 571.070 42.335 585.770 167.400 ;
        RECT 589.670 42.335 604.370 167.400 ;
        RECT 608.270 42.335 638.570 167.400 ;
        RECT 642.470 167.400 694.370 167.640 ;
        RECT 642.470 42.335 657.170 167.400 ;
        RECT 661.070 42.335 675.770 167.400 ;
        RECT 679.670 42.335 694.370 167.400 ;
        RECT 698.270 42.335 728.570 567.820 ;
        RECT 732.470 567.820 818.570 568.060 ;
        RECT 732.470 42.335 747.170 567.820 ;
        RECT 751.070 42.335 765.770 567.820 ;
        RECT 769.670 42.335 784.370 567.820 ;
        RECT 788.270 42.335 818.570 567.820 ;
        RECT 822.470 567.820 908.570 568.060 ;
        RECT 822.470 42.335 837.170 567.820 ;
        RECT 841.070 42.335 855.770 567.820 ;
        RECT 859.670 42.335 874.370 567.820 ;
        RECT 878.270 42.335 908.570 567.820 ;
        RECT 912.470 42.335 927.170 1465.560 ;
        RECT 931.070 42.335 945.770 3355.040 ;
        RECT 949.670 42.335 964.370 3355.040 ;
        RECT 968.270 42.335 998.570 3355.040 ;
        RECT 1002.470 42.335 1017.170 3355.040 ;
        RECT 1021.070 42.335 1035.770 3355.040 ;
        RECT 1039.670 42.335 1054.370 3355.040 ;
        RECT 1058.270 42.335 1088.570 3355.040 ;
        RECT 1092.470 42.335 1107.170 3355.040 ;
        RECT 1111.070 42.335 1125.770 3355.040 ;
        RECT 1129.670 42.335 1144.370 3355.040 ;
        RECT 1148.270 42.335 1178.570 3355.040 ;
        RECT 1182.470 42.335 1197.170 3355.040 ;
        RECT 1201.070 42.335 1215.770 3355.040 ;
        RECT 1219.670 42.335 1234.370 3355.040 ;
        RECT 1238.270 42.335 1268.570 3355.040 ;
        RECT 1272.470 42.335 1287.170 3355.040 ;
        RECT 1291.070 42.335 1305.770 3355.040 ;
        RECT 1309.670 42.335 1324.370 3355.040 ;
        RECT 1328.270 42.335 1358.570 3355.040 ;
        RECT 1362.470 42.335 1377.170 3355.040 ;
        RECT 1381.070 42.335 1395.770 3355.040 ;
        RECT 1399.670 42.335 1414.370 3355.040 ;
        RECT 1418.270 42.335 1448.570 3355.040 ;
        RECT 1452.470 42.335 1467.170 3355.040 ;
        RECT 1471.070 42.335 1485.770 3355.040 ;
        RECT 1489.670 42.335 1504.370 3355.040 ;
        RECT 1508.270 42.335 1538.570 3355.040 ;
        RECT 1542.470 42.335 1557.170 3355.040 ;
        RECT 1561.070 42.335 1575.770 3355.040 ;
        RECT 1579.670 613.220 1594.370 3355.040 ;
        RECT 1598.270 613.220 1628.570 3355.040 ;
        RECT 1579.670 612.980 1628.570 613.220 ;
        RECT 1632.470 613.220 1647.170 3355.040 ;
        RECT 1651.070 613.220 1665.770 3355.040 ;
        RECT 1669.670 613.220 1684.370 3355.040 ;
        RECT 1688.270 3019.580 2205.770 3355.040 ;
        RECT 1688.270 2742.260 1718.570 3019.580 ;
        RECT 1722.470 3019.340 1808.570 3019.580 ;
        RECT 1722.470 2742.500 1737.170 3019.340 ;
        RECT 1741.070 2742.500 1755.770 3019.340 ;
        RECT 1759.670 2742.500 1774.370 3019.340 ;
        RECT 1778.270 2742.500 1808.570 3019.340 ;
        RECT 1722.470 2742.260 1808.570 2742.500 ;
        RECT 1812.470 3019.340 1898.570 3019.580 ;
        RECT 1812.470 2742.500 1827.170 3019.340 ;
        RECT 1831.070 2742.500 1845.770 3019.340 ;
        RECT 1849.670 2742.500 1864.370 3019.340 ;
        RECT 1868.270 2742.500 1898.570 3019.340 ;
        RECT 1812.470 2742.260 1898.570 2742.500 ;
        RECT 1902.470 3019.340 1988.570 3019.580 ;
        RECT 1902.470 2742.500 1917.170 3019.340 ;
        RECT 1921.070 2742.500 1935.770 3019.340 ;
        RECT 1939.670 2742.500 1954.370 3019.340 ;
        RECT 1958.270 2742.500 1988.570 3019.340 ;
        RECT 1902.470 2742.260 1988.570 2742.500 ;
        RECT 1992.470 3019.340 2078.570 3019.580 ;
        RECT 1992.470 2742.500 2007.170 3019.340 ;
        RECT 2011.070 2742.500 2025.770 3019.340 ;
        RECT 2029.670 2742.500 2044.370 3019.340 ;
        RECT 2048.270 2742.500 2078.570 3019.340 ;
        RECT 1992.470 2742.260 2078.570 2742.500 ;
        RECT 2082.470 3019.340 2168.570 3019.580 ;
        RECT 2082.470 2742.500 2097.170 3019.340 ;
        RECT 2101.070 2742.500 2115.770 3019.340 ;
        RECT 2119.670 2742.500 2134.370 3019.340 ;
        RECT 2138.270 2742.500 2168.570 3019.340 ;
        RECT 2082.470 2742.260 2168.570 2742.500 ;
        RECT 2172.470 3019.340 2205.770 3019.580 ;
        RECT 2172.470 2742.500 2187.170 3019.340 ;
        RECT 2191.070 2742.500 2205.770 3019.340 ;
        RECT 2209.670 2742.500 2224.370 3355.040 ;
        RECT 2228.270 2742.500 2258.570 3355.040 ;
        RECT 2172.470 2742.260 2258.570 2742.500 ;
        RECT 2262.470 2742.500 2277.170 3355.040 ;
        RECT 2281.070 2742.500 2295.770 3355.040 ;
        RECT 2299.670 2742.500 2314.370 3355.040 ;
        RECT 2318.270 2742.500 2348.570 3355.040 ;
        RECT 2262.470 2742.260 2348.570 2742.500 ;
        RECT 2352.470 2742.500 2367.170 3355.040 ;
        RECT 2371.070 2742.500 2385.770 3355.040 ;
        RECT 2389.670 2742.500 2404.370 3355.040 ;
        RECT 2408.270 2742.500 2438.570 3355.040 ;
        RECT 2352.470 2742.260 2438.570 2742.500 ;
        RECT 1688.270 2051.320 2438.570 2742.260 ;
        RECT 1688.270 1840.120 1718.570 2051.320 ;
        RECT 1722.470 2051.080 1808.570 2051.320 ;
        RECT 1722.470 1840.360 1737.170 2051.080 ;
        RECT 1741.070 1840.360 1755.770 2051.080 ;
        RECT 1759.670 1840.360 1774.370 2051.080 ;
        RECT 1778.270 1840.360 1808.570 2051.080 ;
        RECT 1722.470 1840.120 1808.570 1840.360 ;
        RECT 1812.470 2051.080 1898.570 2051.320 ;
        RECT 1812.470 1840.360 1827.170 2051.080 ;
        RECT 1831.070 1840.360 1845.770 2051.080 ;
        RECT 1849.670 1840.360 1864.370 2051.080 ;
        RECT 1868.270 1840.360 1898.570 2051.080 ;
        RECT 1812.470 1840.120 1898.570 1840.360 ;
        RECT 1902.470 2051.080 1988.570 2051.320 ;
        RECT 1902.470 1840.360 1917.170 2051.080 ;
        RECT 1921.070 1840.360 1935.770 2051.080 ;
        RECT 1939.670 1840.360 1954.370 2051.080 ;
        RECT 1958.270 1840.360 1988.570 2051.080 ;
        RECT 1902.470 1840.120 1988.570 1840.360 ;
        RECT 1992.470 2051.080 2078.570 2051.320 ;
        RECT 1992.470 1840.360 2007.170 2051.080 ;
        RECT 2011.070 1840.360 2025.770 2051.080 ;
        RECT 2029.670 1840.360 2044.370 2051.080 ;
        RECT 2048.270 1840.360 2078.570 2051.080 ;
        RECT 1992.470 1840.120 2078.570 1840.360 ;
        RECT 2082.470 2051.080 2168.570 2051.320 ;
        RECT 2082.470 1840.360 2097.170 2051.080 ;
        RECT 2101.070 1840.360 2115.770 2051.080 ;
        RECT 2119.670 1840.360 2134.370 2051.080 ;
        RECT 2138.270 1840.360 2168.570 2051.080 ;
        RECT 2082.470 1840.120 2168.570 1840.360 ;
        RECT 2172.470 2051.080 2258.570 2051.320 ;
        RECT 2172.470 1840.360 2187.170 2051.080 ;
        RECT 2191.070 1840.360 2205.770 2051.080 ;
        RECT 2172.470 1840.120 2205.770 1840.360 ;
        RECT 1688.270 1495.300 2205.770 1840.120 ;
        RECT 1688.270 1223.940 1718.570 1495.300 ;
        RECT 1722.470 1495.060 1808.570 1495.300 ;
        RECT 1722.470 1224.180 1737.170 1495.060 ;
        RECT 1741.070 1224.180 1755.770 1495.060 ;
        RECT 1759.670 1224.180 1774.370 1495.060 ;
        RECT 1778.270 1224.180 1808.570 1495.060 ;
        RECT 1722.470 1223.940 1808.570 1224.180 ;
        RECT 1812.470 1495.060 1898.570 1495.300 ;
        RECT 1812.470 1224.180 1827.170 1495.060 ;
        RECT 1831.070 1224.180 1845.770 1495.060 ;
        RECT 1849.670 1224.180 1864.370 1495.060 ;
        RECT 1868.270 1224.180 1898.570 1495.060 ;
        RECT 1812.470 1223.940 1898.570 1224.180 ;
        RECT 1902.470 1495.060 1988.570 1495.300 ;
        RECT 1902.470 1224.180 1917.170 1495.060 ;
        RECT 1921.070 1224.180 1935.770 1495.060 ;
        RECT 1939.670 1224.180 1954.370 1495.060 ;
        RECT 1958.270 1224.180 1988.570 1495.060 ;
        RECT 1902.470 1223.940 1988.570 1224.180 ;
        RECT 1992.470 1495.060 2078.570 1495.300 ;
        RECT 1992.470 1224.180 2007.170 1495.060 ;
        RECT 2011.070 1224.180 2025.770 1495.060 ;
        RECT 2029.670 1224.180 2044.370 1495.060 ;
        RECT 2048.270 1224.180 2078.570 1495.060 ;
        RECT 1992.470 1223.940 2078.570 1224.180 ;
        RECT 2082.470 1495.060 2168.570 1495.300 ;
        RECT 2082.470 1224.180 2097.170 1495.060 ;
        RECT 2101.070 1224.180 2115.770 1495.060 ;
        RECT 2119.670 1224.180 2134.370 1495.060 ;
        RECT 2138.270 1224.180 2168.570 1495.060 ;
        RECT 2082.470 1223.940 2168.570 1224.180 ;
        RECT 2172.470 1495.060 2205.770 1495.300 ;
        RECT 2172.470 1224.180 2187.170 1495.060 ;
        RECT 2191.070 1224.180 2205.770 1495.060 ;
        RECT 2209.670 1224.180 2224.370 2051.080 ;
        RECT 2228.270 1224.180 2258.570 2051.080 ;
        RECT 2172.470 1223.940 2258.570 1224.180 ;
        RECT 2262.470 2051.080 2348.570 2051.320 ;
        RECT 2262.470 1224.180 2277.170 2051.080 ;
        RECT 2281.070 1224.180 2295.770 2051.080 ;
        RECT 2299.670 1224.180 2314.370 2051.080 ;
        RECT 2318.270 1224.180 2348.570 2051.080 ;
        RECT 2262.470 1223.940 2348.570 1224.180 ;
        RECT 2352.470 2051.080 2438.570 2051.320 ;
        RECT 2352.470 1224.180 2367.170 2051.080 ;
        RECT 2371.070 1224.180 2385.770 2051.080 ;
        RECT 2389.670 1224.180 2404.370 2051.080 ;
        RECT 2408.270 1224.180 2438.570 2051.080 ;
        RECT 2352.470 1223.940 2438.570 1224.180 ;
        RECT 1688.270 786.640 2438.570 1223.940 ;
        RECT 1688.270 613.220 1718.570 786.640 ;
        RECT 1632.470 612.980 1718.570 613.220 ;
        RECT 1722.470 786.400 1808.570 786.640 ;
        RECT 1722.470 613.220 1737.170 786.400 ;
        RECT 1741.070 613.220 1755.770 786.400 ;
        RECT 1759.670 613.220 1774.370 786.400 ;
        RECT 1778.270 613.220 1808.570 786.400 ;
        RECT 1722.470 612.980 1808.570 613.220 ;
        RECT 1812.470 786.400 1898.570 786.640 ;
        RECT 1812.470 613.220 1827.170 786.400 ;
        RECT 1831.070 613.220 1845.770 786.400 ;
        RECT 1849.670 613.220 1864.370 786.400 ;
        RECT 1868.270 613.220 1898.570 786.400 ;
        RECT 1812.470 612.980 1898.570 613.220 ;
        RECT 1902.470 786.400 1988.570 786.640 ;
        RECT 1902.470 613.220 1917.170 786.400 ;
        RECT 1921.070 613.220 1935.770 786.400 ;
        RECT 1939.670 613.220 1954.370 786.400 ;
        RECT 1958.270 613.220 1988.570 786.400 ;
        RECT 1902.470 612.980 1988.570 613.220 ;
        RECT 1992.470 786.400 2078.570 786.640 ;
        RECT 1992.470 613.220 2007.170 786.400 ;
        RECT 2011.070 613.220 2025.770 786.400 ;
        RECT 2029.670 613.220 2044.370 786.400 ;
        RECT 2048.270 613.220 2078.570 786.400 ;
        RECT 1992.470 612.980 2078.570 613.220 ;
        RECT 2082.470 786.400 2168.570 786.640 ;
        RECT 2082.470 613.220 2097.170 786.400 ;
        RECT 2101.070 613.220 2115.770 786.400 ;
        RECT 2082.470 612.980 2115.770 613.220 ;
        RECT 1579.670 190.640 2115.770 612.980 ;
        RECT 1579.670 190.400 1628.570 190.640 ;
        RECT 1579.670 42.335 1594.370 190.400 ;
        RECT 1598.270 42.335 1628.570 190.400 ;
        RECT 1632.470 190.400 1718.570 190.640 ;
        RECT 1632.470 42.335 1647.170 190.400 ;
        RECT 1651.070 42.335 1665.770 190.400 ;
        RECT 1669.670 42.335 1684.370 190.400 ;
        RECT 1688.270 42.335 1718.570 190.400 ;
        RECT 1722.470 190.400 1808.570 190.640 ;
        RECT 1722.470 42.335 1737.170 190.400 ;
        RECT 1741.070 42.335 1755.770 190.400 ;
        RECT 1759.670 42.335 1774.370 190.400 ;
        RECT 1778.270 42.335 1808.570 190.400 ;
        RECT 1812.470 190.400 1898.570 190.640 ;
        RECT 1812.470 42.335 1827.170 190.400 ;
        RECT 1831.070 42.335 1845.770 190.400 ;
        RECT 1849.670 42.335 1864.370 190.400 ;
        RECT 1868.270 42.335 1898.570 190.400 ;
        RECT 1902.470 190.400 1988.570 190.640 ;
        RECT 1902.470 42.335 1917.170 190.400 ;
        RECT 1921.070 42.335 1935.770 190.400 ;
        RECT 1939.670 42.335 1954.370 190.400 ;
        RECT 1958.270 42.335 1988.570 190.400 ;
        RECT 1992.470 190.400 2078.570 190.640 ;
        RECT 1992.470 42.335 2007.170 190.400 ;
        RECT 2011.070 42.335 2025.770 190.400 ;
        RECT 2029.670 42.335 2044.370 190.400 ;
        RECT 2048.270 42.335 2078.570 190.400 ;
        RECT 2082.470 190.400 2115.770 190.640 ;
        RECT 2082.470 42.335 2097.170 190.400 ;
        RECT 2101.070 42.335 2115.770 190.400 ;
        RECT 2119.670 42.335 2134.370 786.400 ;
        RECT 2138.270 42.335 2168.570 786.400 ;
        RECT 2172.470 786.400 2258.570 786.640 ;
        RECT 2172.470 42.335 2187.170 786.400 ;
        RECT 2191.070 42.335 2205.770 786.400 ;
        RECT 2209.670 42.335 2224.370 786.400 ;
        RECT 2228.270 42.335 2258.570 786.400 ;
        RECT 2262.470 786.400 2348.570 786.640 ;
        RECT 2262.470 613.220 2277.170 786.400 ;
        RECT 2281.070 613.220 2295.770 786.400 ;
        RECT 2299.670 613.220 2314.370 786.400 ;
        RECT 2318.270 613.220 2348.570 786.400 ;
        RECT 2262.470 612.980 2348.570 613.220 ;
        RECT 2352.470 786.400 2438.570 786.640 ;
        RECT 2352.470 613.220 2367.170 786.400 ;
        RECT 2371.070 613.220 2385.770 786.400 ;
        RECT 2389.670 613.220 2404.370 786.400 ;
        RECT 2408.270 613.220 2438.570 786.400 ;
        RECT 2352.470 612.980 2438.570 613.220 ;
        RECT 2442.470 613.220 2457.170 3355.040 ;
        RECT 2461.070 613.220 2475.770 3355.040 ;
        RECT 2479.670 613.220 2494.370 3355.040 ;
        RECT 2498.270 613.220 2528.570 3355.040 ;
        RECT 2442.470 612.980 2528.570 613.220 ;
        RECT 2532.470 613.220 2547.170 3355.040 ;
        RECT 2551.070 613.220 2565.770 3355.040 ;
        RECT 2569.670 613.220 2584.370 3355.040 ;
        RECT 2588.270 613.220 2618.570 3355.040 ;
        RECT 2532.470 612.980 2618.570 613.220 ;
        RECT 2622.470 613.220 2637.170 3355.040 ;
        RECT 2641.070 613.220 2655.770 3355.040 ;
        RECT 2659.670 613.220 2674.370 3355.040 ;
        RECT 2678.270 613.220 2708.570 3355.040 ;
        RECT 2622.470 612.980 2708.570 613.220 ;
        RECT 2712.470 613.220 2727.170 3355.040 ;
        RECT 2731.070 613.220 2745.770 3355.040 ;
        RECT 2749.670 613.220 2764.370 3355.040 ;
        RECT 2768.270 613.220 2773.160 3355.040 ;
        RECT 2712.470 612.980 2773.160 613.220 ;
        RECT 2262.470 190.640 2773.160 612.980 ;
        RECT 2262.470 190.400 2348.570 190.640 ;
        RECT 2262.470 42.335 2277.170 190.400 ;
        RECT 2281.070 42.335 2295.770 190.400 ;
        RECT 2299.670 42.335 2314.370 190.400 ;
        RECT 2318.270 42.335 2348.570 190.400 ;
        RECT 2352.470 190.400 2438.570 190.640 ;
        RECT 2352.470 42.335 2367.170 190.400 ;
        RECT 2371.070 42.335 2385.770 190.400 ;
        RECT 2389.670 42.335 2404.370 190.400 ;
        RECT 2408.270 42.335 2438.570 190.400 ;
        RECT 2442.470 190.400 2528.570 190.640 ;
        RECT 2442.470 42.335 2457.170 190.400 ;
        RECT 2461.070 42.335 2475.770 190.400 ;
        RECT 2479.670 42.335 2494.370 190.400 ;
        RECT 2498.270 42.335 2528.570 190.400 ;
        RECT 2532.470 190.400 2618.570 190.640 ;
        RECT 2532.470 42.335 2547.170 190.400 ;
        RECT 2551.070 42.335 2565.770 190.400 ;
        RECT 2569.670 42.335 2584.370 190.400 ;
        RECT 2588.270 42.335 2618.570 190.400 ;
        RECT 2622.470 190.400 2708.570 190.640 ;
        RECT 2622.470 42.335 2637.170 190.400 ;
        RECT 2641.070 42.335 2655.770 190.400 ;
        RECT 2659.670 42.335 2674.370 190.400 ;
        RECT 2678.270 42.335 2708.570 190.400 ;
        RECT 2712.470 190.400 2773.160 190.640 ;
        RECT 2712.470 42.335 2727.170 190.400 ;
        RECT 2731.070 42.335 2745.770 190.400 ;
        RECT 2749.670 42.335 2764.370 190.400 ;
        RECT 2768.270 42.335 2773.160 190.400 ;
  END
END user_project_wrapper
END LIBRARY

